* SPICE3 file created from editing.ext - technology: scmos
.include TSMC_180nm.txt

.param SUPPLY=1.8

.option scale=0.09u

M1000 a_2912_n58# ena2c VDD w_2886_n36# CMOSP w=5 l=2
+  ad=55 pd=42 as=8429 ps=5186
M1001 sout0 a_2220_873# a_2100_900# Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=83 ps=64
M1002 a_3163_n518# a_2980_n576# VDD w_3146_n524# CMOSP w=10 l=2
+  ad=210 pd=82 as=0 ps=0
M1003 ena3a a_1092_n417# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=6420 ps=4054
M1004 a_2175_836# a_2131_859# VDD w_2117_852# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1005 enb2a a_1603_n417# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1006 sout3 a_2218_33# a_2098_60# Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=83 ps=64
M1007 a_2218_33# a_2210_n2# gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1008 a_380_n354# s1 gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=54 as=0 ps=0
M1009 a_1748_n4# a_1252_n84# gnd Gnd CMOSN w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1010 a_3711_n46# d2 a_3711_n76# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=168 ps=62
M1011 a_2980_252# enb3c gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1012 gnd a_2175_836# a_2355_831# Gnd CMOSN w=9 l=2
+  ad=0 pd=0 as=63 ps=32
M1013 a_1727_n447# d3 gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1014 a_3304_n443# x3 a_3339_n478# Gnd CMOSN w=10 l=2
+  ad=100 pd=40 as=80 ps=36
M1015 ena2c a_972_n278# VDD w_958_n285# CMOSP w=4 l=2
+  ad=45 pd=38 as=0 ps=0
M1016 d2 a_380_n258# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1017 a_587_n168# a_547_n182# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1018 a_2218_597# a_2210_562# gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1019 x2 a_2900_n58# VDD w_2987_4# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1020 a_1727_n417# b3 a_1727_n447# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1021 sout1 a_2210_562# a_2098_624# w_2221_642# CMOSP w=5 l=2
+  ad=60 pd=44 as=85 ps=64
M1022 a_3661_n330# w3 gnd Gnd CMOSN w=7 l=2
+  ad=126 pd=64 as=0 ps=0
M1023 a_547_n182# d1 a_547_n149# w_529_n155# CMOSP w=9 l=2
+  ad=72 pd=34 as=63 ps=32
M1024 a_3251_495# x3 a_3236_495# Gnd CMOSN w=10 l=2
+  ad=130 pd=46 as=130 ps=46
M1025 a_2980_n576# ena2c gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1026 a_1092_n417# a3 a_1092_n447# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=91 ps=40
M1027 enb1c a_1468_n278# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1028 a_2129_583# ena1as VDD w_2115_576# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1029 a_2126_304# ena2as VDD w_2112_297# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1030 a_2110_60# a_1887_n5# gnd Gnd CMOSN w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1031 a_1603_n417# b2 a_1603_n447# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=91 ps=40
M1032 a_1092_n417# d3 VDD w_1078_n424# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1033 a_2911_n212# ena1c gnd Gnd CMOSN w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1034 a_2882_n382# enb0c VDD w_2885_n338# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1035 ena0as a_693_n145# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1036 a_2975_452# enb0c VDD w_2962_470# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1037 a_2355_831# a_2277_826# gnd Gnd CMOSN w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 a_2353_24# a_2275_n14# VDD w_2335_18# CMOSP w=9 l=2
+  ad=63 pd=32 as=0 ps=0
M1039 a_2980_319# enb2c gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1040 a_1473_n175# a_587_n168# gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1041 a_3221_530# x3 VDD w_3204_524# CMOSP w=10 l=2
+  ad=350 pd=130 as=0 ps=0
M1042 a_2110_624# a_1584_n3# gnd Gnd CMOSN w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1043 a_2881_81# enb3c VDD w_2884_125# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1044 a_3663_329# a_3616_352# VDD w_3602_345# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1045 a_3490_392# x3 VDD w_3473_386# CMOSP w=10 l=2
+  ad=210 pd=82 as=0 ps=0
M1046 a_1326_n145# a_587_n168# VDD w_1312_n152# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1047 VDD b1 a_1464_n417# w_1450_n424# CMOSP w=5 l=2
+  ad=0 pd=0 as=65 ps=36
M1048 a_3065_n592# enb3c VDD w_3051_n599# CMOSP w=5 l=2
+  ad=70 pd=48 as=0 ps=0
M1049 a_2095_345# a_2078_323# a_2107_345# w_2081_367# CMOSP w=5 l=2
+  ad=85 pd=64 as=55 ps=42
M1050 enb3as a_1736_n145# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1051 a_1899_n5# a_1252_n84# VDD w_1873_17# CMOSP w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1052 a_2912_n58# ena2c gnd Gnd CMOSN w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1053 a_3436_n359# a_2975_n443# VDD w_3419_n365# CMOSP w=10 l=2
+  ad=350 pd=130 as=0 ps=0
M1054 a_693_n145# a0 a_693_n175# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=91 ps=40
M1055 a_2275_n14# a_2231_9# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1056 VDD a_2098_60# a_2231_9# w_2217_2# CMOSP w=5 l=2
+  ad=0 pd=0 as=65 ps=36
M1057 a_2207_247# a_2353_555# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1058 a_3490_392# x3 a_3505_357# Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=180 ps=56
M1059 VDD a1 a_826_n278# w_812_n285# CMOSP w=5 l=2
+  ad=0 pd=0 as=65 ps=36
M1060 a_693_n145# a_587_n168# VDD w_679_n152# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1061 a_1435_n1# a_1418_n23# a_1447_n1# w_1421_21# CMOSP w=5 l=2
+  ad=85 pd=64 as=55 ps=42
M1062 a_3634_n79# x1 a_3614_n79# Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=180 ps=56
M1063 and2 a_1843_n566# VDD w_1829_n573# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1064 a_1607_n278# d2 VDD w_1593_n285# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1065 a_3616_352# a_2980_252# VDD w_3602_345# CMOSP w=5 l=2
+  ad=70 pd=48 as=0 ps=0
M1066 ena1as a_831_n145# VDD w_817_n152# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1067 a_3697_480# a_3549_357# a_3682_480# w_3654_474# CMOSP w=7 l=2
+  ad=56 pd=30 as=91 ps=40
M1068 enb0c a_1321_n278# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1069 a_977_n145# a_587_n168# VDD w_963_n152# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1070 VDD b2 a_1607_n278# w_1593_n285# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1071 a_822_n417# d3 VDD w_808_n424# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1072 and1 a_1843_n688# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1073 a_1736_n145# b3 a_1736_n175# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=91 ps=40
M1074 VDD a2 a_977_n145# w_963_n152# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 a_112_n123# s0 VDD w_99_n105# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1076 a_2899_n212# a_2882_n234# ena1c Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=45 ps=38
M1077 a_2098_624# a_2081_602# a_2110_624# w_2084_646# CMOSP w=5 l=2
+  ad=0 pd=0 as=55 ps=42
M1078 a_1887_n5# enb3as a_1252_n84# w_1873_17# CMOSP w=5 l=2
+  ad=85 pd=64 as=120 ps=98
M1079 a_2098_60# a_2081_38# a_1887_n5# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=83 ps=64
M1080 a_2882_n382# enb0c gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1081 a_380_n192# s0 VDD w_366_n199# CMOSP w=5 l=2
+  ad=70 pd=48 as=0 ps=0
M1082 a_1567_n25# enb1as VDD w_1570_19# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1083 a_2247_56# a_2098_60# VDD w_2221_78# CMOSP w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1084 a_2899_n212# a_2882_n234# a_2911_n212# w_2885_n190# CMOSP w=5 l=2
+  ad=60 pd=44 as=55 ps=42
M1085 a_1843_n718# enb1a gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1086 enb1as a_1473_n145# VDD w_1459_n152# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1087 and3 a_1843_n461# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1088 a_1101_n145# a_587_n168# VDD w_1087_n152# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1089 sout0 a_2220_873# a_2249_896# w_2223_918# CMOSP w=5 l=2
+  ad=60 pd=44 as=55 ps=42
M1090 a_2098_60# a_2081_38# a_2110_60# w_2084_82# CMOSP w=5 l=2
+  ad=85 pd=64 as=55 ps=42
M1091 VDD x3 a_3304_n443# w_3287_n449# CMOSP w=10 l=2
+  ad=0 pd=0 as=210 ps=82
M1092 a_2210_562# a_2355_831# VDD w_2337_858# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1093 a_1252_n84# a_1208_n61# VDD w_1194_n68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1094 a_1584_n3# enb1as a_1596_n3# Gnd CMOSN w=5 l=2
+  ad=83 pd=64 as=55 ps=42
M1095 a_972_n308# d2 gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1096 a_2977_n509# ena1c gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1097 w3 a_3163_n518# VDD w_3146_n524# CMOSP w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1098 a_1887_n5# enb3as a_1899_n5# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=55 ps=42
M1099 a_2975_n443# ena0c VDD w_2962_n425# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1100 ena0c a_688_n278# VDD w_674_n285# CMOSP w=4 l=2
+  ad=45 pd=38 as=0 ps=0
M1101 a_1843_n461# ena3a a_1843_n491# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=91 ps=40
M1102 VDD a_1435_n1# a_2131_859# w_2117_852# CMOSP w=5 l=2
+  ad=0 pd=0 as=65 ps=36
M1103 w4 a_3065_n592# VDD w_3051_n599# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1104 a_380_n123# a_112_n178# a_380_n153# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=91 ps=54
M1105 gtr a_3670_450# VDD w_3654_474# CMOSP w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1106 ena0a a_684_n417# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1107 a_2107_345# a_1736_n4# VDD w_2081_367# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1108 a_2900_n58# enb2c ena2c w_2886_n36# CMOSP w=5 l=2
+  ad=60 pd=44 as=0 ps=0
M1109 a_1464_n447# d3 gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1110 a_1096_n308# d2 gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1111 enb0as a_1326_n145# VDD w_1312_n152# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1112 x1 a_2899_n212# VDD w_2986_n150# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1113 a_547_n182# d0 gnd Gnd CMOSN w=9 l=2
+  ad=63 pd=32 as=0 ps=0
M1114 a_1435_n1# enb0as a_1447_n1# Gnd CMOSN w=5 l=2
+  ad=83 pd=64 as=55 ps=42
M1115 a_2975_452# enb0c gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1116 enb3c a_1731_n278# VDD w_1717_n285# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1117 a_831_n145# a_587_n168# VDD w_817_n152# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1118 a_1317_n417# d3 VDD w_1303_n424# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1119 a_2910_103# ena3c gnd Gnd CMOSN w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1120 VDD ena2a a_1843_n566# w_1829_n573# CMOSP w=5 l=2
+  ad=0 pd=0 as=65 ps=36
M1121 a_2095_345# a_2078_323# a_1736_n4# Gnd CMOSN w=5 l=2
+  ad=83 pd=64 as=83 ps=64
M1122 a_1736_n4# enb2as a_1252_n84# w_1722_18# CMOSP w=5 l=2
+  ad=85 pd=64 as=0 ps=0
M1123 a_1719_n26# enb2as VDD w_1722_18# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1124 VDD a_2095_345# a_2228_294# w_2214_287# CMOSP w=5 l=2
+  ad=0 pd=0 as=65 ps=36
M1125 a_3423_395# a_3352_430# gnd Gnd CMOSN w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1126 enb3a a_1727_n417# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1127 VDD a1 a_831_n145# w_817_n152# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 a_2977_386# enb1c VDD w_2964_404# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1129 VDD b0 a_1317_n417# w_1303_n424# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 a_2911_n360# ena0c VDD w_2885_n338# CMOSP w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1131 a_3599_n44# x1 VDD w_3582_n50# CMOSP w=10 l=2
+  ad=210 pd=82 as=0 ps=0
M1132 sout1 a_2210_562# a_2247_620# Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=55 ps=42
M1133 a_3481_n394# x2 a_3466_n394# Gnd CMOSN w=10 l=2
+  ad=120 pd=44 as=130 ps=46
M1134 ena3c a_1096_n278# VDD w_1082_n285# CMOSP w=4 l=2
+  ad=45 pd=38 as=0 ps=0
M1135 a_1612_n145# a_587_n168# VDD w_1598_n152# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1136 a_2126_274# ena2as gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1137 a_3670_480# a_3306_495# VDD w_3654_474# CMOSP w=7 l=2
+  ad=70 pd=34 as=0 ps=0
M1138 a_3490_392# a_2980_319# VDD w_3473_386# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1139 a_684_n417# d3 VDD w_670_n424# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1140 enb2c a_1607_n278# VDD w_1593_n285# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1141 x0 a_2899_n360# VDD w_2986_n298# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1142 VDD a_587_n168# a_1208_n61# w_1194_n68# CMOSP w=5 l=2
+  ad=0 pd=0 as=65 ps=36
M1143 a_3367_395# ena1c a_3352_395# Gnd CMOSN w=10 l=2
+  ad=180 pd=56 as=130 ps=46
M1144 a_3339_n478# x2 a_3319_n478# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=180 ps=56
M1145 a_3616_352# ena3c VDD w_3602_345# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 a_3423_395# a_3352_430# VDD w_3335_424# CMOSP w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1147 ena1a a_822_n417# VDD w_808_n424# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1148 gnd a_2173_n4# a_2353_n9# Gnd CMOSN w=9 l=2
+  ad=0 pd=0 as=63 ps=32
M1149 VDD enb2c a_3163_n518# w_3146_n524# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1150 ena1c a_826_n278# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1151 a_968_n417# d3 VDD w_954_n424# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1152 a_3490_357# a_2980_319# gnd Gnd CMOSN w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1153 a_2129_19# ena3as VDD w_2115_12# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1154 a_3599_n79# x3 gnd Gnd CMOSN w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1155 a_3306_495# a_3221_530# gnd Gnd CMOSN w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1156 gnd d1 a_547_n182# Gnd CMOSN w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1157 a_112_n178# s1 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1158 VDD a2 a_968_n417# w_954_n424# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 a_1843_n795# enb0a VDD w_1829_n802# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1160 d0 a_380_n123# VDD w_366_n130# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1161 a_2249_896# a_2100_900# VDD w_2223_918# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1162 a_2098_624# a_2081_602# a_1584_n3# Gnd CMOSN w=5 l=2
+  ad=83 pd=64 as=0 ps=0
M1163 VDD a_2098_624# a_2231_573# w_2217_566# CMOSP w=5 l=2
+  ad=0 pd=0 as=65 ps=36
M1164 a_2272_271# a_2228_294# VDD w_2214_287# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1165 a_2899_n212# enb1c a_2911_n212# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 VDD ena1c a_3352_430# w_3335_424# CMOSP w=10 l=2
+  ad=0 pd=0 as=210 ps=82
M1167 a_826_n308# d2 gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1168 a_2898_103# a_2881_81# a_2910_103# w_2884_125# CMOSP w=5 l=2
+  ad=60 pd=44 as=55 ps=42
M1169 a_2129_553# ena1as gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1170 enb1a a_1464_n417# VDD w_1450_n424# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1171 a_2112_900# a_1435_n1# gnd Gnd CMOSN w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1172 a_2900_n58# a_2883_n80# ena2c Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=45 ps=38
M1173 a_3306_495# a_3221_530# VDD w_3204_524# CMOSP w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1174 lsr a_3661_n330# VDD w_3645_n306# CMOSP w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1175 ena2a a_968_n417# VDD w_954_n424# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1176 ena2c a_972_n278# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 a_380_n258# a_112_n123# VDD w_366_n265# CMOSP w=5 l=2
+  ad=70 pd=48 as=0 ps=0
M1178 a_3065_n622# a_2980_n643# gnd Gnd CMOSN w=7 l=2
+  ad=133 pd=52 as=0 ps=0
M1179 VDD a0 a_688_n278# w_674_n285# CMOSP w=5 l=2
+  ad=0 pd=0 as=65 ps=36
M1180 a_2244_341# a_2095_345# gnd Gnd CMOSN w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1181 a_2173_n4# a_2129_19# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1182 sout3 a_2210_n2# a_2247_56# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=55 ps=42
M1183 a_2899_n360# enb0c ena0c w_2885_n338# CMOSP w=5 l=2
+  ad=60 pd=44 as=0 ps=0
M1184 a_1736_n4# a_1719_n26# a_1252_n84# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=120 ps=98
M1185 a_1719_n26# enb2as gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1186 a_2210_562# a_2355_831# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1187 a_1473_n145# b1 a_1473_n175# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1188 a_2233_849# a_1252_n84# VDD w_2219_842# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1189 a_2911_n360# ena0c gnd Gnd CMOSN w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1190 a_3673_n300# w2 a_3661_n300# w_3645_n306# CMOSP w=7 l=2
+  ad=91 pd=40 as=70 ps=34
M1191 x3 a_2898_103# VDD w_2985_165# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1192 a_2275_550# a_2231_573# VDD w_2217_566# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1193 a_1731_n278# d2 VDD w_1717_n285# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1194 VDD b0 a_1326_n145# w_1312_n152# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1195 VDD b3 a_1731_n278# w_1717_n285# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1196 a_3661_n330# w4 a_3688_n300# w_3645_n306# CMOSP w=7 l=2
+  ad=63 pd=32 as=56 ps=30
M1197 a_112_n123# s0 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1198 a_2231_9# a_2098_60# a_2231_n21# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=91 ps=40
M1199 VDD enb0c a_3436_n359# w_3419_n365# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1200 a_3616_322# a_2980_252# gnd Gnd CMOSN w=7 l=2
+  ad=133 pd=52 as=0 ps=0
M1201 a_3352_430# x2 a_3387_395# Gnd CMOSN w=10 l=2
+  ad=100 pd=40 as=80 ps=36
M1202 a_2100_900# a_2083_878# a_2112_900# w_2086_922# CMOSP w=5 l=2
+  ad=85 pd=64 as=55 ps=42
M1203 a_2350_276# a_2170_281# a_2350_309# w_2332_303# CMOSP w=9 l=2
+  ad=72 pd=34 as=63 ps=32
M1204 a_3436_n359# x1 VDD w_3419_n365# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1205 a_1843_n596# enb2a gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1206 a_3670_450# a_3549_357# gnd Gnd CMOSN w=7 l=2
+  ad=126 pd=64 as=0 ps=0
M1207 enb0a a_1317_n417# VDD w_1303_n424# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1208 a_2247_620# a_2098_624# gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 VDD a3 a_1096_n278# w_1082_n285# CMOSP w=5 l=2
+  ad=0 pd=0 as=65 ps=36
M1210 a_2173_n4# a_2129_19# VDD w_2115_12# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1211 d3 a_380_n324# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1212 ena3as a_1101_n145# VDD w_1087_n152# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1213 sout2 a_2215_318# a_2244_341# w_2218_363# CMOSP w=5 l=2
+  ad=60 pd=44 as=55 ps=42
M1214 enb2as a_1612_n145# VDD w_1598_n152# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1215 VDD a1 a_822_n417# w_808_n424# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1216 VDD x2 a_3352_430# w_3335_424# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 a_1321_n308# d2 gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1218 a_380_n153# a_112_n123# gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1219 cout a_2353_n9# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1220 a_1603_n417# d3 VDD w_1589_n424# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1221 a_380_n192# a_112_n178# a_380_n222# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=91 ps=54
M1222 a_1447_n1# a_1252_n84# gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1223 a_3221_530# x1 a_3266_495# Gnd CMOSN w=10 l=2
+  ad=90 pd=38 as=120 ps=44
M1224 a_1252_n84# a_1208_n61# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1225 a_1870_n27# enb3as VDD w_1873_17# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1226 a_3304_n443# x2 VDD w_3287_n449# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 a_3163_n518# x3 a_3178_n553# Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=180 ps=56
M1228 a_1321_n278# b0 a_1321_n308# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1229 a_2083_878# ena0as VDD w_2086_922# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1230 a_2081_38# ena3as gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1231 ena2as a_977_n145# VDD w_963_n152# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1232 a_2350_309# a_2272_271# VDD w_2332_303# CMOSP w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1233 a_2899_n360# a_2882_n382# ena0c Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=45 ps=38
M1234 a_1843_n688# ena1a a_1843_n718# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1235 a_3599_n44# x3 VDD w_3582_n50# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1236 a_688_n308# d2 gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1237 a_2175_836# a_2131_859# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1238 and0 a_1843_n795# VDD w_1829_n802# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1239 a_2129_19# a_1887_n5# a_2129_n11# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=91 ps=40
M1240 a_2078_323# ena2as gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1241 a_2215_318# a_2207_247# VDD w_2218_363# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1242 a_3661_n300# w1 VDD w_3645_n306# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1243 a_2975_n443# ena0c gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1244 a_380_n324# s0 VDD w_366_n331# CMOSP w=5 l=2
+  ad=70 pd=48 as=0 ps=0
M1245 d1 a_380_n192# VDD w_366_n199# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1246 a_3221_530# x1 VDD w_3204_524# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1247 a_2210_n2# a_2350_276# VDD w_2332_303# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1248 a_972_n278# a2 a_972_n308# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1249 a_2220_873# a_1252_n84# gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1250 a_2131_859# a_1435_n1# a_2131_829# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=91 ps=40
M1251 a_2898_103# a_2881_81# ena3c Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=45 ps=38
M1252 gtr a_3670_450# gnd Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1253 a_1092_n447# d3 gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1254 a_2272_271# a_2228_294# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1255 sout3 a_2210_n2# a_2098_60# w_2221_78# CMOSP w=5 l=2
+  ad=60 pd=44 as=0 ps=0
M1256 a_2218_33# a_2210_n2# VDD w_2221_78# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1257 a_1584_n3# a_1567_n25# a_1596_n3# w_1570_19# CMOSP w=5 l=2
+  ad=85 pd=64 as=55 ps=42
M1258 a_3549_357# a_3490_392# VDD w_3473_386# CMOSP w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1259 a_2081_602# ena1as gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1260 a_2218_597# a_2210_562# VDD w_2221_642# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1261 VDD a_1736_n4# a_2126_304# w_2112_297# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1262 a_1736_n145# a_587_n168# VDD w_1722_n152# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1263 a_2899_n360# a_2882_n382# a_2911_n360# w_2885_n338# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1264 a_1326_n175# a_587_n168# gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1265 a_1464_n417# b1 a_1464_n447# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1266 ena0c a_688_n278# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1267 a_3549_357# a_3490_392# gnd Gnd CMOSN w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1268 gnd a_2170_281# a_2350_276# Gnd CMOSN w=9 l=2
+  ad=0 pd=0 as=63 ps=32
M1269 a_2228_294# a_2095_345# a_2228_264# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=91 ps=40
M1270 a_1447_n1# a_1252_n84# VDD w_1421_21# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1271 a_3304_n478# a_2977_n509# gnd Gnd CMOSN w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1272 w2 a_3304_n443# gnd Gnd CMOSN w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1273 a_3663_329# a_3616_352# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1274 a_3711_n46# pequ VDD w_3697_n53# CMOSP w=5 l=2
+  ad=70 pd=48 as=0 ps=0
M1275 a_3670_450# a_3306_495# gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1276 a_2110_60# a_1887_n5# VDD w_2084_82# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1277 a_693_n175# a_587_n168# gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1278 sout0 a_1252_n84# a_2100_900# w_2223_918# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1279 a_2275_550# a_2231_573# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1280 a_380_n258# s1 VDD w_366_n265# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1281 cout a_2353_n9# VDD w_2335_18# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1282 VDD a3 a_1101_n145# w_1087_n152# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1283 a_3616_352# ena3c a_3616_322# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1284 VDD b2 a_1612_n145# w_1598_n152# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1285 a_2100_900# a_2083_878# a_1435_n1# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1286 VDD a0 a_684_n417# w_670_n424# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1287 enb3c a_1731_n278# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1288 a_977_n175# a_587_n168# gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1289 a_2131_859# ena0as VDD w_2117_852# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1290 equ a_3711_n46# VDD w_3697_n53# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1291 a_2110_624# a_1584_n3# VDD w_2084_646# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1292 x2 a_2900_n58# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1293 a_822_n447# d3 gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1294 a_2170_281# a_2126_304# VDD w_2112_297# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1295 a_977_n145# a2 a_977_n175# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1296 a_2350_276# a_2272_271# gnd Gnd CMOSN w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1297 a_3065_n592# enb3c a_3065_n622# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1298 a_2231_573# a_2098_624# a_2231_543# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=91 ps=40
M1299 ena3a a_1092_n417# VDD w_1078_n424# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1300 enb2a a_1603_n417# VDD w_1589_n424# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1301 ena3c a_1096_n278# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1302 enb2c a_1607_n278# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1303 a_1468_n278# d2 VDD w_1454_n285# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1304 sout2 a_2215_318# a_2095_345# Gnd CMOSN w=5 l=2
+  ad=58 pd=44 as=0 ps=0
M1305 a_1843_n461# enb3a VDD w_1829_n468# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1306 VDD ena0a a_1843_n795# w_1829_n802# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1307 a_1596_n3# a_1252_n84# gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1308 a_1736_n4# a_1719_n26# a_1748_n4# w_1722_18# CMOSP w=5 l=2
+  ad=0 pd=0 as=55 ps=42
M1309 a_587_n168# a_547_n182# VDD w_529_n155# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1310 VDD b1 a_1468_n278# w_1454_n285# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1311 a_826_n278# a1 a_826_n308# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1312 a_1101_n175# a_587_n168# gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1313 a_2210_n2# a_2350_276# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1314 a_2228_294# a_2207_247# VDD w_2214_287# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1315 a_3436_n359# x3 a_3481_n394# Gnd CMOSN w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1316 a_1607_n308# d2 gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1317 a_2277_826# a_2233_849# VDD w_2219_842# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1318 a_2899_n360# enb0c a_2911_n360# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1319 a_1607_n278# b2 a_1607_n308# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1320 a_2231_9# a_2210_n2# VDD w_2217_2# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1321 a_1899_n5# a_1252_n84# gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1322 a_2980_n576# ena2c VDD w_2967_n558# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1323 a_3670_450# a_3663_329# a_3697_480# w_3654_474# CMOSP w=7 l=2
+  ad=63 pd=32 as=0 ps=0
M1324 a_1208_n61# d1 VDD w_1194_n68# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1325 a_2233_819# a_1252_n84# gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1326 ena0as a_693_n145# VDD w_679_n152# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1327 and2 a_1843_n566# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1328 a_2098_60# ena3as a_1887_n5# w_2084_82# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1329 sout1 a_2218_597# a_2098_624# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1330 a_380_n222# s0 gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1331 ena1as a_831_n145# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1332 a_1584_n3# a_1567_n25# a_1252_n84# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1333 a_3688_n300# w3 a_3673_n300# w_3645_n306# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1334 a_2977_386# enb1c gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1335 a_2231_573# a_2210_562# VDD w_2217_566# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1336 enb3as a_1736_n145# VDD w_1722_n152# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1337 w1 a_3436_n359# gnd Gnd CMOSN w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1338 a_1887_n5# a_1870_n27# a_1252_n84# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1339 a_2980_n643# ena3c VDD w_2967_n625# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1340 a_3711_n46# d2 VDD w_3697_n53# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1341 a_380_n324# s1 VDD w_366_n331# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1342 a_3236_495# ena0c a_3221_495# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=130 ps=46
M1343 a_2900_n58# a_2883_n80# a_2912_n58# w_2886_n36# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1344 a_1727_n417# d3 VDD w_1713_n424# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1345 a_1317_n447# d3 gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1346 a_831_n175# a_587_n168# gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1347 a_2353_555# a_2173_560# a_2353_588# w_2335_582# CMOSP w=9 l=2
+  ad=72 pd=34 as=63 ps=32
M1348 VDD x2 a_3436_n359# w_3419_n365# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1349 a_3304_n443# a_2977_n509# VDD w_3287_n449# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1350 w2 a_3304_n443# VDD w_3287_n449# CMOSP w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1351 a_3163_n553# a_2980_n576# gnd Gnd CMOSN w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1352 enb1as a_1473_n145# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1353 a_2353_n9# a_2173_n4# a_2353_24# w_2335_18# CMOSP w=9 l=2
+  ad=72 pd=34 as=0 ps=0
M1354 a_1843_n566# ena2a a_1843_n596# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1355 a_2881_81# enb3c gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1356 VDD b3 a_1727_n417# w_1713_n424# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1357 a_1317_n417# b0 a_1317_n447# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1358 a_831_n145# a1 a_831_n175# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1359 a_1736_n4# enb2as a_1748_n4# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1360 a_2170_281# a_2126_304# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1361 a_2095_345# ena2as a_2107_345# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=55 ps=42
M1362 a_1612_n175# a_587_n168# gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1363 a_684_n447# d3 gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1364 VDD ena0c a_3221_530# w_3204_524# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1365 a_1208_n61# a_587_n168# a_1208_n91# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=91 ps=40
M1366 VDD a3 a_1092_n417# w_1078_n424# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1367 a_2977_n509# ena1c VDD w_2964_n491# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1368 VDD b2 a_1603_n417# w_1589_n424# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1369 a_2883_n80# enb2c VDD w_2886_n36# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1370 a_2980_319# enb2c VDD w_2967_337# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1371 a_3387_395# x3 a_3367_395# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1372 sout0 a_1252_n84# a_2249_896# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=55 ps=42
M1373 a_968_n447# d3 gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1374 a_2353_588# a_2275_550# VDD w_2335_582# CMOSP w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1375 a_2126_304# a_1736_n4# a_2126_274# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1376 pequ a_3599_n44# gnd Gnd CMOSN w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1377 a_968_n417# a2 a_968_n447# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1378 a_1473_n145# a_587_n168# VDD w_1459_n152# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1379 a_2231_n21# a_2210_n2# gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1380 a_2910_103# ena3c VDD w_2884_125# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1381 VDD ena2c a_3490_392# w_3473_386# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1382 a_2095_345# ena2as a_1736_n4# w_2081_367# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1383 a_3352_430# x3 VDD w_3335_424# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1384 a_2098_624# ena1as a_2110_624# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1385 sout1 a_2218_597# a_2247_620# w_2221_642# CMOSP w=5 l=2
+  ad=0 pd=0 as=55 ps=42
M1386 enb0as a_1326_n145# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1387 x1 a_2899_n212# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1388 a_2207_247# a_2353_555# VDD w_2335_582# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1389 a_3682_480# a_3423_395# a_3670_480# w_3654_474# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1390 a_2353_n9# a_2275_n14# gnd Gnd CMOSN w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1391 a_3505_357# ena2c a_3490_357# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1392 a_2247_56# a_2098_60# gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1393 VDD a0 a_693_n145# w_679_n152# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1394 a_3614_n79# x2 a_3599_n79# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1395 a_1843_n688# enb1a VDD w_1829_n695# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1396 a_380_n258# a_112_n123# a_380_n288# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=91 ps=54
M1397 a_2900_n58# enb2c a_2912_n58# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1398 a_2098_60# ena3as a_2110_60# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1399 a_1887_n5# a_1870_n27# a_1899_n5# w_1873_17# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1400 a_3436_n394# a_2975_n443# gnd Gnd CMOSN w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1401 a_3266_495# x2 a_3251_495# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1402 w4 a_3065_n592# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1403 a_1843_n825# enb0a gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1404 a_2882_n234# enb1c VDD w_2885_n190# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1405 ena0a a_684_n417# VDD w_670_n424# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1406 VDD a_1584_n3# a_2129_583# w_2115_576# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1407 a_2098_624# ena1as a_1584_n3# w_2084_646# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1408 a_972_n278# d2 VDD w_958_n285# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1409 VDD b3 a_1736_n145# w_1722_n152# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1410 a_1326_n145# b0 a_1326_n175# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1411 a_2129_n11# ena3as gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1412 x3 a_2898_103# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1413 ena1a a_822_n417# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1414 a_2275_n14# a_2231_9# VDD w_2217_2# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1415 a_2112_900# a_1435_n1# VDD w_2086_922# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1416 a_3319_n478# enb1c a_3304_n478# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1417 a_2883_n80# enb2c gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1418 lsr a_3661_n330# gnd Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1419 VDD x2 a_3221_530# w_3204_524# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1420 VDD a_2100_900# a_2233_849# w_2219_842# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1421 d0 a_380_n123# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1422 enb3a a_1727_n417# VDD w_1713_n424# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1423 enb1c a_1468_n278# VDD w_1454_n285# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1424 a_688_n278# a0 a_688_n308# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1425 a_2131_829# ena0as gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1426 a_2107_345# a_1736_n4# gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1427 a_2244_341# a_2095_345# VDD w_2218_363# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1428 sout3 a_2218_33# a_2247_56# w_2221_78# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1429 a_1096_n278# d2 VDD w_1082_n285# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1430 enb1a a_1464_n417# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1431 gnd w2 a_3661_n330# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1432 a_3163_n518# x3 VDD w_3146_n524# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1433 x0 a_2899_n360# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1434 a_822_n417# a1 a_822_n447# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1435 ena2a a_968_n417# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1436 a_2173_560# a_2129_583# VDD w_2115_576# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1437 a_1731_n308# d2 gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1438 d2 a_380_n258# VDD w_366_n265# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1439 a_2249_896# a_2100_900# gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1440 gnd a_2173_560# a_2353_555# Gnd CMOSN w=9 l=2
+  ad=0 pd=0 as=63 ps=32
M1441 a_1418_n23# enb0as gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1442 a_1603_n447# d3 gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1443 a_1435_n1# enb0as a_1252_n84# w_1421_21# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1444 a_1418_n23# enb0as VDD w_1421_21# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1445 a_1731_n278# b3 a_1731_n308# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1446 gnd w4 a_3661_n330# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1447 a_112_n178# s1 VDD w_99_n160# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1448 a_2228_264# a_2207_247# gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1449 VDD ena3a a_1843_n461# w_1829_n468# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1450 a_3599_n44# x0 a_3634_n79# Gnd CMOSN w=10 l=2
+  ad=100 pd=40 as=0 ps=0
M1451 a_380_n123# a_112_n178# VDD w_366_n130# CMOSP w=5 l=2
+  ad=70 pd=48 as=0 ps=0
M1452 w3 a_3163_n518# gnd Gnd CMOSN w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1453 pequ a_3599_n44# VDD w_3582_n50# CMOSP w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1454 a_2247_620# a_2098_624# VDD w_2221_642# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1455 gnd a_3663_329# a_3670_450# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1456 a_1096_n278# a3 a_1096_n308# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1457 a_1464_n417# d3 VDD w_1450_n424# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1458 a_380_n324# s0 a_380_n354# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1459 a_1435_n1# a_1418_n23# a_1252_n84# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1460 enb0c a_1321_n278# VDD w_1307_n285# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1461 a_2353_555# a_2275_550# gnd Gnd CMOSN w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1462 a_3352_395# a_2977_386# gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1463 a_1596_n3# a_1252_n84# VDD w_1570_19# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1464 and1 a_1843_n688# VDD w_1829_n695# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1465 VDD x2 a_3599_n44# w_3582_n50# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1466 a_826_n278# d2 VDD w_812_n285# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1467 enb0a a_1317_n417# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1468 a_2081_38# ena3as VDD w_2084_82# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1469 a_2355_831# a_2175_836# a_2355_864# w_2337_858# CMOSP w=9 l=2
+  ad=72 pd=34 as=63 ps=32
M1470 a_2898_103# enb3c a_2910_103# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1471 a_2980_252# enb3c VDD w_2967_270# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1472 a_2231_543# a_2210_562# gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1473 a_1567_n25# enb1as gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1474 a_2980_n643# ena3c gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1475 ena3as a_1101_n145# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1476 enb2as a_1612_n145# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1477 a_3352_430# a_2977_386# VDD w_3335_424# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1478 a_2078_323# ena2as VDD w_2081_367# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1479 a_2882_n234# enb1c gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1480 a_1736_n175# a_587_n168# gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1481 VDD a_1887_n5# a_2129_19# w_2115_12# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1482 a_3661_n330# w1 gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1483 a_3065_n592# a_2980_n643# VDD w_3051_n599# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1484 a_1870_n27# enb3as gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1485 ena2as a_977_n145# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1486 VDD enb1c a_3304_n443# w_3287_n449# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1487 a_3178_n553# enb2c a_3163_n553# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1488 a_3711_n76# pequ gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1489 a_2898_103# enb3c ena3c w_2884_125# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1490 a_1584_n3# enb1as a_1252_n84# w_1570_19# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1491 a_2355_864# a_2277_826# VDD w_2337_858# CMOSP w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1492 a_380_n288# s1 gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1493 d3 a_380_n324# VDD w_366_n331# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1494 a_1101_n145# a3 a_1101_n175# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1495 a_1612_n145# b2 a_1612_n175# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1496 a_684_n417# a0 a_684_n447# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1497 a_2911_n212# ena1c VDD w_2885_n190# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1498 a_2100_900# ena0as a_2112_900# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1499 a_2081_602# ena1as VDD w_2084_646# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1500 and3 a_1843_n461# VDD w_1829_n468# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1501 a_1748_n4# a_1252_n84# VDD w_1722_18# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1502 VDD b1 a_1473_n145# w_1459_n152# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1503 a_3436_n359# x3 VDD w_3419_n365# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1504 a_1843_n491# enb3a gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1505 sout2 a_2207_247# a_2244_341# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1506 a_3221_495# a_2975_452# gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1507 a_2220_873# a_1252_n84# VDD w_2223_918# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1508 gnd a_3423_395# a_3670_450# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1509 and0 a_1843_n795# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1510 VDD x0 a_3599_n44# w_3582_n50# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1511 a_1321_n278# d2 VDD w_1307_n285# CMOSP w=5 l=2
+  ad=65 pd=36 as=0 ps=0
M1512 a_2173_560# a_2129_583# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1513 a_380_n192# a_112_n178# VDD w_366_n199# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1514 d1 a_380_n192# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1515 VDD b0 a_1321_n278# w_1307_n285# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1516 a_2100_900# ena0as a_1435_n1# w_2086_922# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1517 a_2083_878# ena0as gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1518 VDD ena1a a_1843_n688# w_1829_n695# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1519 a_688_n278# d2 VDD w_674_n285# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1520 a_3221_530# a_2975_452# VDD w_3204_524# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1521 a_2277_826# a_2233_849# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1522 a_1843_n566# enb2a VDD w_1829_n573# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1523 a_1208_n91# d1 gnd Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1524 a_3451_n394# enb0c a_3436_n394# Gnd CMOSN w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1525 a_2215_318# a_2207_247# gnd Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1526 a_2129_583# a_1584_n3# a_2129_553# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1527 ena1c a_826_n278# VDD w_812_n285# CMOSP w=4 l=2
+  ad=45 pd=38 as=0 ps=0
M1528 a_1468_n308# d2 gnd Gnd CMOSN w=7 l=2
+  ad=91 pd=40 as=0 ps=0
M1529 a_547_n149# d0 VDD w_529_n155# CMOSP w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1530 sout2 a_2207_247# a_2095_345# w_2218_363# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1531 a_3466_n394# x1 a_3451_n394# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1532 a_1843_n795# ena0a a_1843_n825# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1533 w1 a_3436_n359# VDD w_3419_n365# CMOSP w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1534 a_1468_n278# b1 a_1468_n308# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1535 equ a_3711_n46# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1536 VDD a2 a_972_n278# w_958_n285# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1537 a_2899_n212# enb1c ena1c w_2885_n190# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1538 a_2233_849# a_2100_900# a_2233_819# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1539 a_380_n123# a_112_n123# VDD w_366_n130# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
C0 ena3c a_2980_n643# 0.01fF
C1 a_1870_n27# a_1252_n84# 0.14fF
C2 VDD a_2231_573# 0.03fF
C3 a_1870_n27# VDD 0.03fF
C4 w_3051_n599# a_3065_n592# 0.14fF
C5 x2 a_2980_252# 0.07fF
C6 w_3146_n524# a_3163_n518# 0.11fF
C7 enb1as w_1459_n152# 0.03fF
C8 a_2126_304# VDD 0.03fF
C9 gnd ena2a 0.24fF
C10 w_2967_n558# a_2980_n576# 0.03fF
C11 x2 enb0c 0.06fF
C12 w_2086_922# a_2100_900# 0.13fF
C13 w_1829_n695# VDD 0.22fF
C14 w_3654_474# a_3663_329# 0.06fF
C15 w_2221_642# a_2210_562# 0.16fF
C16 a_587_n168# b0 0.10fF
C17 w_1722_18# a_1736_n4# 0.13fF
C18 enb3c a_2881_81# 0.32fF
C19 enb2c a_2883_n80# 0.32fF
C20 ena1c a_2911_n212# 0.28fF
C21 x3 a_2975_n443# 0.01fF
C22 w_2117_852# gnd 0.09fF
C23 w_3419_n365# a_2975_n443# 0.06fF
C24 w_3645_n306# w1 0.06fF
C25 a_2277_826# w_2219_842# 0.03fF
C26 a_2275_n14# VDD 0.07fF
C27 w_2086_922# VDD 0.08fF
C28 a_1584_n3# a_2110_624# 0.28fF
C29 w_2337_858# a_2277_826# 0.11fF
C30 a_2231_9# VDD 0.03fF
C31 a_2228_294# a_2207_247# 0.04fF
C32 enb1c a_3304_n443# 0.08fF
C33 w_2081_367# a_2107_345# 0.07fF
C34 w_812_n285# a1 0.07fF
C35 w_2214_287# a_2095_345# 0.07fF
C36 x3 a_2980_319# 0.07fF
C37 s0 s1 0.56fF
C38 d1 a_547_n182# 0.20fF
C39 a_112_n178# a_380_n123# 0.43fF
C40 gnd ena1a 0.26fF
C41 w_3287_n449# a_3304_n443# 0.11fF
C42 gnd enb2as 0.10fF
C43 a_3221_530# a_3306_495# 0.03fF
C44 a_2350_276# a_2170_281# 0.20fF
C45 a_2975_452# enb0c 0.02fF
C46 a_2218_33# w_2221_78# 0.12fF
C47 a_2173_n4# w_2335_18# 0.06fF
C48 b1 a_1468_n278# 0.10fF
C49 x0 a_3599_n44# 0.08fF
C50 w_3146_n524# VDD 0.30fF
C51 w_366_n130# VDD 0.23fF
C52 enb0c a_2899_n360# 0.08fF
C53 a_2098_624# a_2231_573# 0.10fF
C54 b2 ena3c 0.01fF
C55 w_3582_n50# x0 0.06fF
C56 VDD a_2980_n643# 0.07fF
C57 sout0 a_2249_896# 0.70fF
C58 ena2c ena3c 12.26fF
C59 gnd x1 0.50fF
C60 a_1435_n1# a_1418_n23# 0.08fF
C61 w_1717_n285# enb3c 0.03fF
C62 ena2as d1 0.01fF
C63 a_2081_602# VDD 0.03fF
C64 a_1887_n5# ena3as 1.26fF
C65 a_2247_56# gnd 0.28fF
C66 a_2098_60# a_2210_n2# 0.23fF
C67 w4 a_3661_n330# 0.08fF
C68 a_2899_n360# a_2911_n360# 0.70fF
C69 a_1899_n5# enb3as 0.25fF
C70 a_3423_395# a_3490_392# 0.01fF
C71 a_2112_900# a_2100_900# 0.70fF
C72 w_2967_337# gnd 0.01fF
C73 gnd w3 0.14fF
C74 a_2277_826# gnd 0.16fF
C75 cout gnd 0.04fF
C76 VDD w_2967_270# 0.10fF
C77 gnd a_684_n417# 0.03fF
C78 a_2100_900# a_2233_849# 0.10fF
C79 a_1887_n5# a_2098_60# 1.27fF
C80 x2 a_3221_530# 0.08fF
C81 w_2115_576# ena1as 0.09fF
C82 VDD ena3c 0.44fF
C83 a1 a_826_n278# 0.10fF
C84 a_1887_n5# a_1899_n5# 0.70fF
C85 VDD a_1208_n61# 0.03fF
C86 a_2175_836# a_1252_n84# 0.00fF
C87 a_2175_836# VDD 0.07fF
C88 b2 ena2c 0.01fF
C89 gnd a_3670_450# 0.11fF
C90 a_2112_900# VDD 0.06fF
C91 VDD a_3163_n518# 0.03fF
C92 gnd a_1101_n145# 0.03fF
C93 gnd ena0c 0.31fF
C94 w_529_n155# a_587_n168# 0.03fF
C95 VDD a_1727_n417# 0.03fF
C96 d2 b0 0.11fF
C97 a_1252_n84# a_2233_849# 0.04fF
C98 VDD a_2233_849# 0.03fF
C99 b2 a_1603_n417# 0.10fF
C100 gnd a_2882_n382# 0.16fF
C101 b0 a_1321_n278# 0.10fF
C102 VDD w_1087_n152# 0.22fF
C103 a_2083_878# gnd 0.04fF
C104 gnd enb3c 0.21fF
C105 a_2081_602# w_2084_646# 0.12fF
C106 x3 x2 2.48fF
C107 ena0c x1 0.07fF
C108 w_1194_n68# d1 0.10fF
C109 VDD b2 0.17fF
C110 a_2098_624# a_2081_602# 0.08fF
C111 w_3419_n365# x2 0.06fF
C112 VDD ena2c 0.35fF
C113 a_1252_n84# a_2100_900# 0.23fF
C114 VDD a_2100_900# 0.59fF
C115 a_2977_n509# a_3163_n518# 0.01fF
C116 a_1736_n4# a_1748_n4# 0.70fF
C117 w_1598_n152# a_1612_n145# 0.10fF
C118 enb2as a_587_n168# 0.00fF
C119 w_2084_82# a_1887_n5# 0.22fF
C120 gnd and0 0.04fF
C121 x3 w2 0.01fF
C122 gnd a_587_n168# 0.10fF
C123 w_1303_n424# enb0a 0.03fF
C124 b2 d3 0.11fF
C125 gnd a_3423_395# 0.06fF
C126 ena1c ena3c 0.06fF
C127 w_99_n160# gnd 0.08fF
C128 gnd a_380_n222# 0.34fF
C129 VDD a_1603_n417# 0.03fF
C130 b3 a_1736_n145# 0.10fF
C131 gnd s1 0.20fF
C132 a_2170_281# w_2112_297# 0.03fF
C133 w_2962_470# VDD 0.11fF
C134 a_1252_n84# VDD 1.14fF
C135 a_1567_n25# gnd 0.04fF
C136 gnd a_2882_n234# 0.16fF
C137 gnd enb2c 0.43fF
C138 gnd a_2249_896# 0.28fF
C139 a_2098_60# w_2221_78# 0.22fF
C140 w_817_n152# VDD 0.22fF
C141 a_1584_n3# gnd 0.08fF
C142 VDD d3 0.76fF
C143 d2 w_1717_n285# 0.10fF
C144 ena0a a_1843_n795# 0.10fF
C145 w_2081_367# a_1736_n4# 0.22fF
C146 gnd and1 0.04fF
C147 ena2c a_2900_n58# 1.32fF
C148 ena3c a_2898_103# 1.32fF
C149 ena0c a_2882_n382# 0.14fF
C150 w_2115_576# a_2173_560# 0.03fF
C151 w_2115_12# VDD 0.22fF
C152 ena2as a_2095_345# 0.08fF
C153 b2 ena1c 0.01fF
C154 gnd and2 0.04fF
C155 ena1c ena2c 13.78fF
C156 w_2217_566# a_2231_573# 0.10fF
C157 ena0c enb3c 0.08fF
C158 sout1 a_2247_620# 0.70fF
C159 a_380_n324# a_380_n354# 0.15fF
C160 VDD a_2977_n509# 0.08fF
C161 w_1450_n424# enb1a 0.03fF
C162 w_2885_n338# ena0c 0.22fF
C163 w_1829_n802# VDD 0.22fF
C164 a_1447_n1# w_1421_21# 0.07fF
C165 a1 a_831_n145# 0.10fF
C166 b3 enb0c 0.01fF
C167 a_2170_281# a_2272_271# 0.28fF
C168 w_2967_337# enb2c 0.06fF
C169 w_1312_n152# a_587_n168# 0.10fF
C170 w_954_n424# VDD 0.22fF
C171 w_2886_n36# enb2c 0.16fF
C172 a_3423_395# a_3670_450# 0.08fF
C173 gnd a_2107_345# 0.28fF
C174 a_1596_n3# a_1252_n84# 0.28fF
C175 a_1596_n3# VDD 0.06fF
C176 x2 a_2977_386# 0.01fF
C177 x3 a_3352_430# 0.08fF
C178 a_1418_n23# gnd 0.04fF
C179 a_2207_247# VDD 0.35fF
C180 w_2885_n338# a_2882_n382# 0.12fF
C181 gnd enb1c 0.72fF
C182 VDD a_2900_n58# 0.16fF
C183 w_1598_n152# enb2as 0.03fF
C184 w_366_n130# d0 0.03fF
C185 w_954_n424# d3 0.10fF
C186 VDD ena1c 0.30fF
C187 a_1736_n4# a_2078_323# 0.14fF
C188 w_2084_646# VDD 0.08fF
C189 a_2098_624# VDD 0.59fF
C190 a_2355_831# a_2210_562# 0.02fF
C191 w_1593_n285# enb2c 0.03fF
C192 gnd and3 0.04fF
C193 ena0c enb2c 0.21fF
C194 w_1087_n152# a3 0.07fF
C195 gnd w_2335_18# 0.21fF
C196 VDD a_1464_n417# 0.03fF
C197 d2 gnd 0.20fF
C198 w_1713_n424# b3 0.07fF
C199 ena1as a_2110_624# 0.25fF
C200 a_1435_n1# ena1as 0.05fF
C201 a3 ena2c 0.01fF
C202 w_808_n424# VDD 0.22fF
C203 w_1713_n424# enb3a 0.03fF
C204 enb2c enb3c 0.11fF
C205 a_1719_n26# enb2as 0.30fF
C206 w_366_n331# VDD 0.27fF
C207 gnd equ 0.04fF
C208 w_958_n285# a2 0.07fF
C209 a_112_n123# a_112_n178# 0.14fF
C210 gnd a_1719_n26# 0.04fF
C211 w_2335_582# a_2275_550# 0.11fF
C212 gnd a_1321_n278# 0.03fF
C213 a_2228_294# a_2095_345# 0.10fF
C214 VDD a_2898_103# 0.16fF
C215 a_2210_562# a_2247_620# 0.24fF
C216 w_99_n160# s1 0.06fF
C217 VDD a_688_n278# 0.03fF
C218 w4 a_3065_n592# 0.02fF
C219 w_674_n285# VDD 0.22fF
C220 w_808_n424# d3 0.10fF
C221 w_366_n331# d3 0.03fF
C222 w_3697_n53# a_3711_n46# 0.14fF
C223 cout w_2335_18# 0.03fF
C224 w_3645_n306# VDD 0.19fF
C225 s0 a_380_n324# 0.28fF
C226 w_2962_n425# VDD 0.11fF
C227 VDD a3 0.17fF
C228 w_2218_363# VDD 0.08fF
C229 ena0c enb1c 0.08fF
C230 a_2173_560# w_2335_582# 0.06fF
C231 VDD a_2975_n443# 0.34fF
C232 VDD ena3a 0.07fF
C233 a_2110_60# gnd 0.28fF
C234 a3 d3 0.11fF
C235 a_2899_n212# a_2911_n212# 0.70fF
C236 w_679_n152# ena0as 0.03fF
C237 a_2098_624# w_2084_646# 0.13fF
C238 w_3602_345# a_3616_352# 0.14fF
C239 w_2884_125# ena3c 0.22fF
C240 enb1c enb3c 0.14fF
C241 a_2129_19# gnd 0.03fF
C242 gnd a_3599_n44# 0.03fF
C243 a_2173_n4# a_2210_n2# 0.00fF
C244 a_1584_n3# a_1567_n25# 0.08fF
C245 gnd a_1096_n278# 0.03fF
C246 VDD a_2980_319# 0.07fF
C247 w_1593_n285# d2 0.10fF
C248 a_2081_38# gnd 0.04fF
C249 VDD d1 0.31fF
C250 a_2350_276# gnd 0.12fF
C251 x1 a_3599_n44# 0.08fF
C252 gnd a_2980_n576# 0.25fF
C253 w_2218_363# a_2207_247# 0.16fF
C254 w_1598_n152# a_587_n168# 0.10fF
C255 x2 ena3c 0.06fF
C256 w_2964_404# gnd 0.01fF
C257 gnd a_977_n145# 0.03fF
C258 a_2098_60# a_2231_9# 0.10fF
C259 a_2173_n4# a_2353_n9# 0.20fF
C260 VDD d0 0.16fF
C261 a_2173_560# a_2210_562# 0.00fF
C262 w_3582_n50# x1 0.06fF
C263 a_2218_33# VDD 0.03fF
C264 VDD a_968_n417# 0.03fF
C265 a_1435_n1# a_1447_n1# 0.70fF
C266 VDD a_1473_n145# 0.03fF
C267 a3 ena1c 0.01fF
C268 enb0as a_1252_n84# 0.09fF
C269 VDD a_693_n145# 0.03fF
C270 enb0as VDD 0.16fF
C271 enb1c a_2882_n234# 0.32fF
C272 w_99_n105# a_112_n123# 0.03fF
C273 enb1c enb2c 11.82fF
C274 gnd a_3616_352# 0.06fF
C275 a_2215_318# VDD 0.03fF
C276 gnd a_972_n278# 0.03fF
C277 w_3335_424# x3 0.06fF
C278 sout1 a_2218_597# 0.08fF
C279 w_2337_858# a_2355_831# 0.09fF
C280 VDD a_3306_495# 0.17fF
C281 a_1736_n4# enb2as 0.08fF
C282 w_1829_n695# a_1843_n688# 0.10fF
C283 a_1736_n4# gnd 0.08fF
C284 a_1317_n417# enb0a 0.02fF
C285 x3 x0 0.07fF
C286 a_2220_873# a_2100_900# 0.14fF
C287 VDD w_2217_566# 0.22fF
C288 ena1c a_2980_319# 0.08fF
C289 w_1589_n424# b2 0.07fF
C290 w_2332_303# VDD 0.22fF
C291 w_674_n285# a_688_n278# 0.10fF
C292 x2 ena2c 0.06fF
C293 VDD a_3661_n330# 0.04fF
C294 w_954_n424# a_968_n417# 0.10fF
C295 w_2884_125# VDD 0.09fF
C296 VDD a_822_n417# 0.03fF
C297 w_3473_386# a_3490_392# 0.11fF
C298 gnd a_380_n123# 0.01fF
C299 gnd b1 0.31fF
C300 enb0c a_3436_n359# 0.08fF
C301 w_2115_576# a_2129_583# 0.10fF
C302 w_1589_n424# a_1603_n417# 0.10fF
C303 gnd a0 0.32fF
C304 gnd a_2912_n58# 0.28fF
C305 w_1722_n152# b3 0.07fF
C306 a_2215_318# a_2207_247# 0.16fF
C307 w_2885_n190# a_2911_n212# 0.07fF
C308 a_2220_873# a_1252_n84# 0.16fF
C309 gnd a_380_n324# 0.01fF
C310 w_2962_n425# a_2975_n443# 0.03fF
C311 a_2220_873# VDD 0.03fF
C312 w_3051_n599# enb3c 0.07fF
C313 ena1as gnd 0.05fF
C314 w_1570_19# a_1567_n25# 0.12fF
C315 w_1589_n424# VDD 0.22fF
C316 w_3287_n449# enb1c 0.06fF
C317 VDD x2 0.19fF
C318 w_1454_n285# VDD 0.22fF
C319 a_2355_831# gnd 0.01fF
C320 ena3as w_1087_n152# 0.03fF
C321 a_2218_33# sout3 0.08fF
C322 w_963_n152# a_587_n168# 0.10fF
C323 w_3204_524# a_3221_530# 0.13fF
C324 w_1570_19# a_1584_n3# 0.13fF
C325 ena2a enb0a 0.01fF
C326 w_1589_n424# d3 0.10fF
C327 w_1307_n285# b0 0.07fF
C328 w_366_n265# s1 0.07fF
C329 w_2886_n36# a_2912_n58# 0.07fF
C330 a_2218_597# a_2210_562# 0.16fF
C331 a0 a_684_n417# 0.10fF
C332 enb1as a_1252_n84# 0.09fF
C333 x2 a_2977_n509# 0.01fF
C334 x3 a_3304_n443# 0.08fF
C335 w_3602_345# a_2980_252# 0.07fF
C336 enb1as VDD 0.16fF
C337 a_2098_624# w_2217_566# 0.07fF
C338 gnd a_2910_103# 0.28fF
C339 gnd a_1736_n145# 0.03fF
C340 gnd w_2112_297# 0.09fF
C341 w_3335_424# a_2977_386# 0.06fF
C342 gnd a_2247_620# 0.28fF
C343 a_2353_555# w_2335_582# 0.09fF
C344 w_366_n130# a_112_n178# 0.12fF
C345 gnd a_826_n278# 0.03fF
C346 VDD a_3663_329# 0.07fF
C347 ena3as a_1252_n84# 0.09fF
C348 ena3as VDD 0.19fF
C349 w_2985_165# x3 0.03fF
C350 b0 a_1326_n145# 0.10fF
C351 VDD a_2095_345# 0.59fF
C352 w_2962_470# a_2975_452# 0.03fF
C353 VDD a_2975_452# 0.27fF
C354 b1 ena0c 0.01fF
C355 enb2c a_2980_n576# 0.20fF
C356 w_3204_524# x3 0.06fF
C357 ena1a enb0a 0.01fF
C358 w_2218_363# a_2215_318# 0.12fF
C359 w_2081_367# ena2as 0.16fF
C360 gnd enb0a 0.17fF
C361 x2 ena1c 0.19fF
C362 VDD a_2899_n360# 0.16fF
C363 a_2098_60# VDD 0.59fF
C364 VDD a_1731_n278# 0.03fF
C365 w_808_n424# a_822_n417# 0.10fF
C366 w_2115_12# ena3as 0.09fF
C367 a_1899_n5# a_1252_n84# 0.28fF
C368 w_2884_125# a_2898_103# 0.13fF
C369 a_2131_859# VDD 0.03fF
C370 a_1899_n5# VDD 0.06fF
C371 b2 a_1607_n278# 0.10fF
C372 enb1as a_1596_n3# 0.25fF
C373 gnd a_2980_252# 0.25fF
C374 gnd a_2275_550# 0.16fF
C375 s0 a_112_n123# 0.13fF
C376 d1 d0 0.30fF
C377 VDD a_1843_n795# 0.03fF
C378 w_3645_n306# a_3661_n330# 0.09fF
C379 gnd a_1447_n1# 0.28fF
C380 gnd enb0c 0.54fF
C381 gnd a_2272_271# 0.16fF
C382 a_1435_n1# ena2as 0.06fF
C383 a_587_n168# b1 0.10fF
C384 w_1082_n285# ena3c 0.03fF
C385 VDD a_380_n192# 0.11fF
C386 a_2207_247# a_2095_345# 0.23fF
C387 a_2244_341# VDD 0.06fF
C388 a_587_n168# a0 0.10fF
C389 gnd enb3as 0.11fF
C390 a_2210_n2# gnd 0.86fF
C391 ena2as a_2078_323# 0.30fF
C392 gnd a_2911_n360# 0.28fF
C393 VDD a2 0.17fF
C394 gnd a_2173_560# 0.35fF
C395 w_2964_404# enb1c 0.06fF
C396 x1 a_2980_252# 0.07fF
C397 ena1as a_587_n168# 0.01fF
C398 x1 enb0c 0.16fF
C399 gnd a_1092_n417# 0.03fF
C400 VDD a_2899_n212# 0.16fF
C401 s1 a_380_n324# 0.05fF
C402 w_1829_n468# VDD 0.22fF
C403 VDD a_1607_n278# 0.03fF
C404 a_1887_n5# gnd 0.08fF
C405 w_3654_474# a_3670_450# 0.09fF
C406 w_366_n265# d2 0.03fF
C407 a2 d3 0.11fF
C408 pequ a_3711_n46# 0.05fF
C409 w_1829_n802# a_1843_n795# 0.10fF
C410 w_2217_2# a_2210_n2# 0.09fF
C411 enb2c a_2912_n58# 0.25fF
C412 w_2084_82# VDD 0.08fF
C413 x2 a_2975_n443# 0.01fF
C414 enb3c a_2910_103# 0.25fF
C415 x3 a_3436_n359# 0.08fF
C416 a_2247_56# a_2210_n2# 0.24fF
C417 a_2353_n9# gnd 0.10fF
C418 w_3419_n365# a_3436_n359# 0.13fF
C419 VDD a_1843_n688# 0.03fF
C420 w_3645_n306# w2 0.06fF
C421 a_1736_n4# a_2107_345# 0.28fF
C422 w_2986_n298# VDD 0.08fF
C423 VDD a_1843_n566# 0.03fF
C424 a_1584_n3# ena1as 1.22fF
C425 b3 ena3c 0.01fF
C426 w_1873_17# enb3as 0.16fF
C427 w1 a_3436_n359# 0.03fF
C428 w_1722_18# a_1252_n84# 0.22fF
C429 w_2967_n558# ena2c 0.06fF
C430 w_2967_n625# a_2980_n643# 0.03fF
C431 w_2964_n491# gnd 0.01fF
C432 w_1722_18# VDD 0.08fF
C433 a_2244_341# a_2207_247# 0.24fF
C434 a_2098_60# sout3 1.20fF
C435 w_954_n424# a2 0.07fF
C436 ena0c a_2980_252# 0.07fF
C437 ena1c a_3352_430# 0.08fF
C438 a_2210_562# a_2231_573# 0.04fF
C439 x2 a_2980_319# 0.07fF
C440 x3 a_3490_392# 0.08fF
C441 VDD a1 0.17fF
C442 gnd a_831_n145# 0.03fF
C443 ena0c enb0c 0.01fF
C444 a_380_n258# a_380_n288# 0.15fF
C445 a_2275_n14# a_2173_n4# 0.28fF
C446 VDD a_112_n178# 0.30fF
C447 VDD w_1829_n573# 0.22fF
C448 b3 a_1727_n417# 0.10fF
C449 w_1873_17# a_1887_n5# 0.13fF
C450 VDD a_1468_n278# 0.03fF
C451 w_1459_n152# a_587_n168# 0.10fF
C452 w_817_n152# a1 0.07fF
C453 w_2218_363# a_2095_345# 0.22fF
C454 w_3654_474# a_3423_395# 0.06fF
C455 a1 d3 0.11fF
C456 a2 ena1c 0.01fF
C457 w_679_n152# a_587_n168# 0.10fF
C458 a_1727_n417# enb3a 0.02fF
C459 enb0c a_2882_n382# 0.34fF
C460 w_1082_n285# VDD 0.22fF
C461 ena0c a_2911_n360# 0.28fF
C462 ena1c a_2899_n212# 1.32fF
C463 w_2967_n625# ena3c 0.06fF
C464 w_2223_918# a_2100_900# 0.22fF
C465 w_2967_n558# VDD 0.10fF
C466 w_3582_n50# a_3599_n44# 0.11fF
C467 enb0c enb3c 0.13fF
C468 VDD a_3065_n592# 0.16fF
C469 w_529_n155# a_547_n182# 0.09fF
C470 w_2221_642# a_2247_620# 0.07fF
C471 gnd a_3221_530# 0.05fF
C472 VDD a_1843_n461# 0.03fF
C473 w_2885_n338# enb0c 0.16fF
C474 VDD w_1303_n424# 0.22fF
C475 b3 ena2c 0.01fF
C476 w_2115_576# VDD 0.22fF
C477 gnd a_1326_n145# 0.03fF
C478 a_1736_n4# a_1719_n26# 0.08fF
C479 d2 w_812_n285# 0.10fF
C480 a_3549_357# a_3490_392# 0.03fF
C481 d2 b1 0.11fF
C482 w_366_n199# VDD 0.31fF
C483 w_963_n152# a_977_n145# 0.10fF
C484 w_2086_922# ena0as 0.16fF
C485 gnd w4 0.20fF
C486 w_1829_n695# enb1a 0.10fF
C487 d2 a0 0.11fF
C488 w_1303_n424# d3 0.10fF
C489 w_2885_n338# a_2911_n360# 0.07fF
C490 x1 a_3221_530# 0.08fF
C491 gnd ena0a 0.22fF
C492 w_2223_918# a_1252_n84# 0.16fF
C493 VDD a_3711_n46# 0.12fF
C494 w_2223_918# VDD 0.08fF
C495 ena3as d1 0.01fF
C496 a_2218_597# gnd 0.22fF
C497 gnd a_112_n123# 0.04fF
C498 a_1435_n1# w_2086_922# 0.22fF
C499 w_2218_363# a_2244_341# 0.07fF
C500 w_2885_n190# VDD 0.09fF
C501 a_1252_n84# w_1421_21# 0.22fF
C502 VDD w_1421_21# 0.08fF
C503 VDD b3 0.17fF
C504 a_2170_281# VDD 0.07fF
C505 gnd a_547_n182# 0.01fF
C506 w_2986_n150# VDD 0.08fF
C507 enb0c enb2c 0.15fF
C508 gnd x3 1.15fF
C509 w_670_n424# a_684_n417# 0.10fF
C510 VDD enb3a 0.07fF
C511 b3 d3 0.11fF
C512 w3 w4 0.01fF
C513 w_3335_424# VDD 0.28fF
C514 w2 a_3661_n330# 0.08fF
C515 a_2215_318# a_2095_345# 0.14fF
C516 a_2218_33# a_2098_60# 0.14fF
C517 a_3670_450# gtr 0.05fF
C518 a_2247_56# w_2221_78# 0.07fF
C519 w_1829_n468# ena3a 0.07fF
C520 w_99_n105# VDD 0.08fF
C521 a_684_n417# ena0a 0.02fF
C522 gnd w1 0.06fF
C523 w_808_n424# a1 0.07fF
C524 gnd ena2as 0.05fF
C525 ena0c a_3221_530# 0.08fF
C526 x3 x1 0.30fF
C527 VDD w_2967_n625# 0.09fF
C528 VDD x0 0.07fF
C529 w_2987_4# VDD 0.11fF
C530 w_3419_n365# x1 0.06fF
C531 w_1312_n152# a_1326_n145# 0.10fF
C532 x2 w2 0.10fF
C533 x3 w3 0.21fF
C534 a_1603_n417# enb2a 0.02fF
C535 gnd a_2353_555# 0.08fF
C536 a_2207_247# a_2170_281# 0.00fF
C537 gnd a_3549_357# 0.06fF
C538 enb0c enb1c 12.75fF
C539 gnd a_380_n258# 0.01fF
C540 VDD enb2a 0.07fF
C541 a_1748_n4# a_1252_n84# 0.28fF
C542 w_2885_n190# ena1c 0.22fF
C543 a_2112_900# ena0as 0.25fF
C544 a_1748_n4# VDD 0.06fF
C545 a2 a_968_n417# 0.10fF
C546 b3 ena1c 0.01fF
C547 w_2335_582# VDD 0.18fF
C548 w_1082_n285# a3 0.07fF
C549 w_1450_n424# b1 0.07fF
C550 gnd a_2911_n212# 0.28fF
C551 b0 ena3c 0.01fF
C552 a_1435_n1# a_2112_900# 0.28fF
C553 ena0c x3 0.10fF
C554 w_3335_424# ena1c 0.06fF
C555 w_2987_4# a_2900_n58# 0.06fF
C556 gnd a_2129_583# 0.03fF
C557 a_2173_n4# VDD 0.07fF
C558 ena2c a_2883_n80# 0.14fF
C559 ena3c a_2881_81# 0.14fF
C560 ena3a a_1843_n461# 0.10fF
C561 ena0as a_2100_900# 0.08fF
C562 gnd a_2977_386# 0.36fF
C563 gnd a_2228_294# 0.03fF
C564 a_1435_n1# a_2100_900# 1.27fF
C565 sout1 a_2098_624# 1.20fF
C566 a_587_n168# a_547_n182# 0.02fF
C567 gnd a_1870_n27# 0.04fF
C568 w_2081_367# VDD 0.08fF
C569 gnd a_2231_573# 0.03fF
C570 a_3549_357# a_3670_450# 0.08fF
C571 w_2985_165# VDD 0.08fF
C572 a_2126_304# gnd 0.03fF
C573 VDD a_2210_562# 0.32fF
C574 a_2173_n4# w_2115_12# 0.03fF
C575 a_2353_n9# w_2335_18# 0.09fF
C576 w_2335_582# a_2207_247# 0.03fF
C577 x1 a_2977_386# 0.01fF
C578 x2 a_3352_430# 0.08fF
C579 w_1829_n695# ena1a 0.07fF
C580 x3 a_3423_395# 0.01fF
C581 b0 ena2c 0.01fF
C582 VDD w_3204_524# 0.30fF
C583 ena0as VDD 0.19fF
C584 VDD a_2883_n80# 0.06fF
C585 w_2221_642# a_2218_597# 0.12fF
C586 w_366_n199# d1 0.03fF
C587 ena2as a_587_n168# 0.01fF
C588 a_1435_n1# a_1252_n84# 1.31fF
C589 a_2098_60# ena3as 0.08fF
C590 a_2110_624# VDD 0.06fF
C591 a_1435_n1# VDD 0.27fF
C592 ena3a enb3a 0.10fF
C593 a_2275_n14# gnd 0.16fF
C594 sout0 a_2100_900# 1.20fF
C595 a_2078_323# VDD 0.03fF
C596 VDD enb1a 0.07fF
C597 VDD b0 0.17fF
C598 a_2231_9# gnd 0.03fF
C599 a1 a_822_n417# 0.10fF
C600 w_1873_17# a_1870_n27# 0.12fF
C601 a_1736_n4# w_2112_297# 0.07fF
C602 a_1887_n5# a_2110_60# 0.28fF
C603 w_1307_n285# d2 0.10fF
C604 a_2207_247# a_2210_562# 0.13fF
C605 ena0c a_2977_386# 0.01fF
C606 w_2217_2# a_2275_n14# 0.03fF
C607 b0 d3 0.10fF
C608 w_3602_345# ena3c 0.07fF
C609 d2 w_3697_n53# 0.10fF
C610 a_1584_n3# ena2as 0.07fF
C611 a_1887_n5# a_2129_19# 0.10fF
C612 a_2244_341# a_2095_345# 0.28fF
C613 VDD s0 0.10fF
C614 VDD a_2881_81# 0.06fF
C615 a_2350_276# a_2210_n2# 0.02fF
C616 sout0 a_1252_n84# 0.08fF
C617 w_812_n285# a_826_n278# 0.10fF
C618 s1 a_380_n258# 0.05fF
C619 w_2217_2# a_2231_9# 0.10fF
C620 b2 a_1612_n145# 0.10fF
C621 w_1722_n152# a_587_n168# 0.10fF
C622 w_1307_n285# a_1321_n278# 0.10fF
C623 w_2337_858# a_2175_836# 0.06fF
C624 w_2219_842# a_2233_849# 0.10fF
C625 w_3697_n53# equ 0.03fF
C626 a_2900_n58# a_2883_n80# 0.08fF
C627 a_2081_38# a_1887_n5# 0.14fF
C628 enb0as w_1421_21# 0.16fF
C629 w_1078_n424# a_1092_n417# 0.10fF
C630 gnd a_2980_n643# 0.25fF
C631 a_2098_624# a_2210_562# 0.23fF
C632 ena3a enb2a 0.01fF
C633 ena2c a_3490_392# 0.08fF
C634 gnd a_2081_602# 0.04fF
C635 w_1459_n152# b1 0.07fF
C636 x3 enb1c 0.07fF
C637 VDD a_3436_n359# 0.03fF
C638 w_1454_n285# a_1468_n278# 0.10fF
C639 w_2117_852# a_2175_836# 0.03fF
C640 VDD a_1317_n417# 0.03fF
C641 w_2084_82# ena3as 0.16fF
C642 w_3287_n449# x3 0.06fF
C643 ena2as a_2107_345# 0.25fF
C644 a_2100_900# w_2219_842# 0.07fF
C645 w_679_n152# a0 0.07fF
C646 w_2084_646# a_2110_624# 0.07fF
C647 w_1194_n68# a_587_n168# 0.07fF
C648 gnd w_2967_270# 0.01fF
C649 a_2098_624# a_2110_624# 0.70fF
C650 VDD a_1612_n145# 0.03fF
C651 w_2332_303# a_2170_281# 0.06fF
C652 b0 ena1c 0.01fF
C653 w_3146_n524# w3 0.02fF
C654 w_2985_165# a_2898_103# 0.06fF
C655 gnd ena3c 0.29fF
C656 VDD a_3490_392# 0.03fF
C657 w_2084_82# a_2098_60# 0.13fF
C658 gnd a_1208_n61# 0.03fF
C659 b1 enb0c 0.01fF
C660 w_2223_918# a_2220_873# 0.12fF
C661 w_1717_n285# VDD 0.22fF
C662 w_2986_n298# a_2899_n360# 0.06fF
C663 a_2175_836# gnd 0.35fF
C664 a_1252_n84# w_2219_842# 0.09fF
C665 a_1584_n3# a_2129_583# 0.10fF
C666 gnd a_2112_900# 0.28fF
C667 gnd a_380_n153# 0.34fF
C668 gnd a_3163_n518# 0.03fF
C669 a_1464_n417# enb1a 0.02fF
C670 VDD w_2219_842# 0.22fF
C671 x1 ena3c 0.06fF
C672 gnd a_1727_n417# 0.03fF
C673 a_2083_878# w_2086_922# 0.12fF
C674 gnd a_2233_849# 0.03fF
C675 VDD ena2a 0.07fF
C676 w_2337_858# VDD 0.18fF
C677 w_3602_345# VDD 0.23fF
C678 w_529_n155# VDD 0.18fF
C679 d2 w_958_n285# 0.10fF
C680 enb1c a_2911_n212# 0.25fF
C681 w_3051_n599# w4 0.03fF
C682 w_2117_852# VDD 0.22fF
C683 gnd b2 0.31fF
C684 gnd ena2c 0.26fF
C685 gnd a_2100_900# 0.16fF
C686 w_3335_424# x2 0.06fF
C687 a_2277_826# a_2175_836# 0.28fF
C688 w_366_n331# s0 0.28fF
C689 d2 a_380_n258# 0.02fF
C690 w_366_n265# a_112_n123# 0.28fF
C691 w3 a_3163_n518# 0.03fF
C692 a_2898_103# a_2881_81# 0.08fF
C693 w_1829_n695# and1 0.03fF
C694 ena3a enb1a 0.01fF
C695 x2 x0 0.07fF
C696 a_112_n178# a_380_n192# 0.28fF
C697 w_2987_4# x2 0.03fF
C698 ena0as d1 0.01fF
C699 ena0c ena3c 0.07fF
C700 gnd a_1603_n417# 0.03fF
C701 x1 ena2c 0.06fF
C702 w_3582_n50# x3 0.06fF
C703 enb2as a_1252_n84# 0.14fF
C704 w_954_n424# ena2a 0.03fF
C705 enb2as VDD 0.15fF
C706 VDD ena1a 0.07fF
C707 gnd a_1252_n84# 1.27fF
C708 gnd VDD 6.54fF
C709 w_2967_270# enb3c 0.06fF
C710 w_2886_n36# ena2c 0.22fF
C711 w_1589_n424# enb2a 0.03fF
C712 ena2as w_963_n152# 0.03fF
C713 ena3c enb3c 0.14fF
C714 gnd d3 0.19fF
C715 w_3146_n524# enb2c 0.06fF
C716 b3 a_1731_n278# 0.10fF
C717 VDD x1 0.20fF
C718 w_2217_2# VDD 0.22fF
C719 w_366_n199# a_380_n192# 0.13fF
C720 gnd w_2115_12# 0.09fF
C721 w_1087_n152# a_1101_n145# 0.10fF
C722 w_1829_n573# a_1843_n566# 0.10fF
C723 a_1435_n1# enb0as 0.08fF
C724 a_2247_56# VDD 0.06fF
C725 w_3204_524# a_3306_495# 0.02fF
C726 w_1593_n285# b2 0.07fF
C727 w_1829_n468# a_1843_n461# 0.10fF
C728 gnd a_2977_n509# 0.36fF
C729 a_2210_562# w_2217_566# 0.09fF
C730 w_670_n424# a0 0.07fF
C731 w_2214_287# a_2272_271# 0.03fF
C732 b2 ena0c 0.01fF
C733 a_587_n168# a_1208_n61# 0.10fF
C734 ena0c ena2c 0.13fF
C735 w_2886_n36# VDD 0.09fF
C736 a_1584_n3# a_2081_602# 0.14fF
C737 w_2967_337# VDD 0.10fF
C738 a_2277_826# VDD 0.07fF
C739 cout VDD 0.07fF
C740 w_366_n265# a_380_n258# 0.13fF
C741 w_1873_17# a_1252_n84# 0.22fF
C742 VDD a_684_n417# 0.03fF
C743 w_1873_17# VDD 0.08fF
C744 a_112_n123# a_380_n123# 0.05fF
C745 a_2173_560# a_2275_550# 0.28fF
C746 gnd a_1596_n3# 0.28fF
C747 gnd a_2207_247# 1.98fF
C748 a_2275_n14# w_2335_18# 0.11fF
C749 enb0c a_2911_n360# 0.25fF
C750 x2 a_3304_n443# 0.08fF
C751 ena3c enb2c 0.07fF
C752 gnd a_2900_n58# 0.11fF
C753 ena2c enb3c 0.08fF
C754 w_3335_424# a_3352_430# 0.11fF
C755 a_2083_878# a_2100_900# 0.08fF
C756 w_3645_n306# lsr 0.02fF
C757 w_2885_n190# a_2899_n212# 0.13fF
C758 gnd ena1c 0.20fF
C759 w_2986_n150# a_2899_n212# 0.06fF
C760 w_1593_n285# VDD 0.22fF
C761 VDD a_3670_450# 0.04fF
C762 w_1312_n152# VDD 0.22fF
C763 VDD a_1101_n145# 0.03fF
C764 w_1087_n152# a_587_n168# 0.10fF
C765 w2 a_3304_n443# 0.03fF
C766 w_958_n285# a_972_n278# 0.10fF
C767 VDD ena0c 0.43fF
C768 a_2098_624# gnd 0.16fF
C769 a_1736_n4# ena2as 1.23fF
C770 enb2c a_3163_n518# 0.08fF
C771 w_3204_524# x2 0.06fF
C772 a_1887_n5# enb3as 0.08fF
C773 a_587_n168# b2 0.10fF
C774 w_1829_n468# enb3a 0.10fF
C775 ena2c a_3423_395# 0.01fF
C776 gnd a_1464_n417# 0.03fF
C777 ena0c d3 4.36fF
C778 x1 ena1c 0.01fF
C779 w_366_n199# a_112_n178# 0.28fF
C780 VDD a_2882_n382# 0.05fF
C781 VDD enb3c 0.15fF
C782 a_2083_878# VDD 0.03fF
C783 w_808_n424# ena1a 0.03fF
C784 w_3654_474# gtr 0.02fF
C785 w_2886_n36# a_2900_n58# 0.13fF
C786 w_2885_n338# VDD 0.09fF
C787 w_2884_125# a_2881_81# 0.12fF
C788 w_2964_404# a_2977_386# 0.03fF
C789 gnd a_2898_103# 0.11fF
C790 ena3c enb1c 0.02fF
C791 ena2c enb2c 0.20fF
C792 VDD and0 0.07fF
C793 a_2100_900# a_2249_896# 0.28fF
C794 VDD a_587_n168# 0.81fF
C795 sout3 a_2247_56# 0.70fF
C796 w_2081_367# a_2095_345# 0.13fF
C797 gnd a_688_n278# 0.03fF
C798 VDD a_3423_395# 0.09fF
C799 w_1307_n285# enb0c 0.03fF
C800 w_99_n160# VDD 0.10fF
C801 w_2962_n425# gnd 0.01fF
C802 gnd a3 0.31fF
C803 w_529_n155# d1 0.06fF
C804 w_2986_n298# x0 0.03fF
C805 w_817_n152# a_587_n168# 0.10fF
C806 w_3204_524# a_2975_452# 0.06fF
C807 sout0 a_2220_873# 0.08fF
C808 gnd a_2975_n443# 0.19fF
C809 ena0a enb0a 0.19fF
C810 ena0c ena1c 14.33fF
C811 w_529_n155# d0 0.11fF
C812 gnd ena3a 0.24fF
C813 a_1567_n25# a_1252_n84# 0.14fF
C814 a_1567_n25# VDD 0.03fF
C815 VDD a_2882_n234# 0.05fF
C816 a_1435_n1# ena3as 0.09fF
C817 VDD enb2c 0.28fF
C818 a_1252_n84# a_2249_896# 0.24fF
C819 VDD a_2249_896# 0.06fF
C820 a_1584_n3# a_1252_n84# 1.38fF
C821 a_1584_n3# VDD 0.29fF
C822 w_3473_386# x3 0.06fF
C823 w_1829_n802# and0 0.03fF
C824 w_2221_642# VDD 0.08fF
C825 x2 a_3436_n359# 0.08fF
C826 x1 a_2975_n443# 0.14fF
C827 ena2as w_2112_297# 0.09fF
C828 a_2078_323# a_2095_345# 0.08fF
C829 b2 enb1c 0.01fF
C830 gnd a_2980_319# 0.54fF
C831 ena2c enb1c 0.01fF
C832 ena1c enb3c 0.04fF
C833 a_2131_859# ena0as 0.04fF
C834 w_1722_18# a_1748_n4# 0.07fF
C835 VDD and1 0.07fF
C836 w_1598_n152# b2 0.07fF
C837 w_3645_n306# w3 0.06fF
C838 a_2126_304# a_1736_n4# 0.10fF
C839 VDD and2 0.07fF
C840 gnd d1 0.18fF
C841 a_3661_n330# lsr 0.05fF
C842 a_1435_n1# a_2131_859# 0.10fF
C843 ena1as a_2129_583# 0.04fF
C844 enb2c a_2977_n509# 0.01fF
C845 w_1829_n573# enb2a 0.10fF
C846 x3 a_2980_252# 0.07fF
C847 gnd d0 0.07fF
C848 x1 a_2980_319# 0.07fF
C849 w_3051_n599# a_2980_n643# 0.07fF
C850 a_2218_33# gnd 0.22fF
C851 a_2107_345# VDD 0.06fF
C852 w_3146_n524# a_2980_n576# 0.06fF
C853 gnd a_968_n417# 0.03fF
C854 w_2221_78# a_2210_n2# 0.16fF
C855 gnd a_1473_n145# 0.03fF
C856 x3 enb0c 0.06fF
C857 w_674_n285# ena0c 0.03fF
C858 a_1418_n23# a_1252_n84# 0.14fF
C859 a_1418_n23# VDD 0.03fF
C860 d2 b2 0.11fF
C861 gnd a_693_n145# 0.03fF
C862 w_3419_n365# enb0c 0.06fF
C863 VDD enb1c 0.42fF
C864 enb0as gnd 0.04fF
C865 w_3473_386# a_3549_357# 0.02fF
C866 w_2962_n425# ena0c 0.06fF
C867 a3 a_1101_n145# 0.10fF
C868 a3 ena0c 0.01fF
C869 w_3654_474# a_3549_357# 0.06fF
C870 w_2967_337# a_2980_319# 0.03fF
C871 w_1722_n152# a_1736_n145# 0.10fF
C872 w_1598_n152# VDD 0.22fF
C873 a_3599_n44# pequ 0.03fF
C874 a_1584_n3# a_1596_n3# 0.70fF
C875 gnd a_2215_318# 0.22fF
C876 ena1c a_2882_n234# 0.14fF
C877 enb3c a_2898_103# 0.08fF
C878 enb2c a_2900_n58# 0.08fF
C879 w_3287_n449# VDD 0.31fF
C880 w_3582_n50# pequ 0.02fF
C881 ena1c enb2c 0.18fF
C882 gnd a_3306_495# 0.06fF
C883 VDD and3 0.07fF
C884 w_2335_18# VDD 0.18fF
C885 a_1584_n3# w_2084_646# 0.22fF
C886 a_1584_n3# a_2098_624# 1.27fF
C887 enb1c a_2977_n509# 0.09fF
C888 w_2221_642# a_2098_624# 0.22fF
C889 d2 VDD 0.96fF
C890 w_2332_303# gnd 0.24fF
C891 w_366_n331# s1 0.07fF
C892 s0 a_380_n192# 0.05fF
C893 gnd a_3661_n330# 0.11fF
C894 ena0c a_2980_319# 0.07fF
C895 gnd a_822_n417# 0.03fF
C896 w_3287_n449# a_2977_n509# 0.06fF
C897 VDD equ 0.07fF
C898 a_587_n168# a3 0.10fF
C899 a_1719_n26# a_1252_n84# 0.14fF
C900 a_1719_n26# VDD 0.03fF
C901 VDD a_1321_n278# 0.03fF
C902 a_2353_555# a_2173_560# 0.20fF
C903 a_2126_304# w_2112_297# 0.10fF
C904 w_366_n130# a_380_n123# 0.13fF
C905 w_1570_19# a_1252_n84# 0.22fF
C906 ena3c a_3616_352# 0.08fF
C907 w_3602_345# a_3663_329# 0.03fF
C908 w_1570_19# VDD 0.08fF
C909 gnd a_2220_873# 0.22fF
C910 w_1722_n152# enb3as 0.03fF
C911 ena1c enb1c 0.14fF
C912 w_1717_n285# a_1731_n278# 0.10fF
C913 w_670_n424# ena0a 0.03fF
C914 w_1312_n152# enb0as 0.03fF
C915 gnd x2 0.69fF
C916 w3 a_3661_n330# 0.08fF
C917 a_3423_395# a_2980_319# 0.01fF
C918 a_2110_60# VDD 0.06fF
C919 ena2c a_2980_n576# 0.02fF
C920 sout2 a_2207_247# 0.08fF
C921 gnd w2 0.15fF
C922 ena1as a_2081_602# 0.30fF
C923 d1 a_587_n168# 0.16fF
C924 w_2214_287# a_2228_294# 0.10fF
C925 x2 x1 0.86fF
C926 a_2129_19# VDD 0.03fF
C927 x3 a_3221_530# 0.08fF
C928 VDD w_963_n152# 0.22fF
C929 VDD a_1096_n278# 0.03fF
C930 b1 ena3c 0.01fF
C931 w_366_n265# VDD 0.26fF
C932 w_3582_n50# VDD 0.31fF
C933 w_3051_n599# VDD 0.26fF
C934 gnd enb1as 0.11fF
C935 a_2081_38# VDD 0.03fF
C936 a_1870_n27# enb3as 0.30fF
C937 w_1570_19# a_1596_n3# 0.07fF
C938 gnd a_3663_329# 0.10fF
C939 w_1303_n424# b0 0.07fF
C940 a_380_n123# a_380_n153# 0.15fF
C941 w_2117_852# a_2131_859# 0.10fF
C942 enb0as a_587_n168# 0.01fF
C943 VDD a_2980_n576# 0.08fF
C944 gnd a_2095_345# 0.16fF
C945 gnd ena3as 0.05fF
C946 gnd a_2975_452# 0.23fF
C947 a_2129_19# w_2115_12# 0.10fF
C948 w_2964_404# VDD 0.10fF
C949 w_1078_n424# VDD 0.22fF
C950 VDD a_977_n145# 0.03fF
C951 a_1435_n1# w_1421_21# 0.13fF
C952 w_1450_n424# VDD 0.22fF
C953 a_1887_n5# a_1870_n27# 0.08fF
C954 gnd a_2899_n360# 0.11fF
C955 w_2884_125# enb3c 0.16fF
C956 a_2098_60# gnd 0.16fF
C957 w_1078_n424# d3 0.10fF
C958 a_2355_831# a_2175_836# 0.20fF
C959 gnd a_1731_n278# 0.03fF
C960 ena0c x2 0.11fF
C961 w_366_n199# s0 0.07fF
C962 VDD a_3616_352# 0.16fF
C963 w_3419_n365# x3 0.06fF
C964 w_674_n285# d2 0.10fF
C965 gnd a_2131_859# 0.03fF
C966 a_2977_n509# a_2980_n576# 0.01fF
C967 w_1450_n424# d3 0.10fF
C968 a_1899_n5# gnd 0.28fF
C969 VDD a_972_n278# 0.03fF
C970 sout1 a_2210_562# 0.08fF
C971 b1 ena2c 0.01fF
C972 w_2218_363# sout2 0.13fF
C973 w_2223_918# sout0 0.13fF
C974 d2 a3 0.11fF
C975 gnd a_1843_n795# 0.03fF
C976 ena3c a_2910_103# 0.28fF
C977 ena2a a_1843_n566# 0.10fF
C978 ena2c a_2912_n58# 0.28fF
C979 a_1736_n4# a_1252_n84# 1.39fF
C980 a_2231_9# a_2210_n2# 0.04fF
C981 w_1303_n424# a_1317_n417# 0.10fF
C982 w_2217_2# a_2098_60# 0.07fF
C983 gnd a_3352_430# 0.03fF
C984 a_1736_n4# VDD 0.29fF
C985 w_3419_n365# w1 0.02fF
C986 a_2098_60# a_2247_56# 0.28fF
C987 gnd a_380_n192# 0.01fF
C988 a_2244_341# gnd 0.28fF
C989 a_112_n123# a_380_n258# 0.28fF
C990 gnd a2 0.31fF
C991 VDD a_380_n123# 0.11fF
C992 VDD w_812_n285# 0.22fF
C993 w_1829_n573# ena2a 0.07fF
C994 a_3663_329# a_3670_450# 0.08fF
C995 VDD b1 0.17fF
C996 gnd a_2899_n212# 0.11fF
C997 a_1418_n23# enb0as 0.30fF
C998 gnd a_1607_n278# 0.03fF
C999 VDD a0 0.15fF
C1000 VDD a_2912_n58# 0.06fF
C1001 w_99_n105# s0 0.06fF
C1002 w_1873_17# a_1899_n5# 0.07fF
C1003 w_2967_270# a_2980_252# 0.03fF
C1004 ena1as a_1252_n84# 0.06fF
C1005 VDD a_380_n324# 0.11fF
C1006 ena1as VDD 0.19fF
C1007 b1 d3 0.11fF
C1008 ena1a a_1843_n688# 0.10fF
C1009 a0 d3 0.11fF
C1010 gnd a_1843_n688# 0.03fF
C1011 ena0c a_2899_n360# 1.32fF
C1012 gnd a_1843_n566# 0.03fF
C1013 w_817_n152# ena1as 0.03fF
C1014 enb0c ena3c 10.54fF
C1015 a_380_n324# d3 0.02fF
C1016 w_1722_18# enb2as 0.16fF
C1017 enb1as a_587_n168# 0.01fF
C1018 w_1450_n424# a_1464_n417# 0.10fF
C1019 a3 a_1096_n278# 0.10fF
C1020 a_2899_n360# a_2882_n382# 0.08fF
C1021 w_3473_386# ena2c 0.06fF
C1022 w_1717_n285# b3 0.07fF
C1023 gnd a1 0.31fF
C1024 ena3as a_587_n168# 0.01fF
C1025 gnd a_112_n178# 0.04fF
C1026 sout2 a_2215_318# 0.08fF
C1027 x3 a_2977_386# 0.01fF
C1028 w_2885_n338# a_2899_n360# 0.13fF
C1029 gnd a_1468_n278# 0.03fF
C1030 VDD a_2910_103# 0.06fF
C1031 a_1567_n25# enb1as 0.30fF
C1032 VDD a_1736_n145# 0.03fF
C1033 w_812_n285# ena1c 0.03fF
C1034 VDD w_2112_297# 0.22fF
C1035 VDD a_2247_620# 0.06fF
C1036 w_1078_n424# a3 0.07fF
C1037 b1 ena1c 0.01fF
C1038 VDD a_826_n278# 0.03fF
C1039 a2 ena0c 0.01fF
C1040 gnd w_2967_n558# 0.01fF
C1041 a_1584_n3# enb1as 0.08fF
C1042 a_2900_n58# a_2912_n58# 0.70fF
C1043 gnd a_3065_n592# 0.05fF
C1044 w_1078_n424# ena3a 0.03fF
C1045 ena2c a_2980_252# 0.10fF
C1046 w_1593_n285# a_1607_n278# 0.10fF
C1047 VDD w_1459_n152# 0.22fF
C1048 w_3654_474# VDD 0.19fF
C1049 b2 enb0c 0.01fF
C1050 gnd a_1843_n461# 0.03fF
C1051 w_3473_386# VDD 0.24fF
C1052 x2 enb1c 0.07fF
C1053 enb0c ena2c 0.04fF
C1054 a_1435_n1# ena0as 1.29fF
C1055 w_2081_367# a_2078_323# 0.12fF
C1056 a_1584_n3# ena3as 0.10fF
C1057 w_1454_n285# enb1c 0.03fF
C1058 w_679_n152# VDD 0.22fF
C1059 w_2115_576# gnd 0.09fF
C1060 b1 a_1464_n417# 0.10fF
C1061 VDD enb0a 0.07fF
C1062 ena1as w_2084_646# 0.16fF
C1063 w_3287_n449# x2 0.06fF
C1064 a_2098_624# ena1as 0.08fF
C1065 a_2126_304# ena2as 0.04fF
C1066 a_3352_430# a_3423_395# 0.03fF
C1067 gnd a_3711_n46# 0.01fF
C1068 w_1713_n424# a_1727_n417# 0.10fF
C1069 w_3287_n449# w2 0.02fF
C1070 a_380_n192# a_380_n222# 0.15fF
C1071 VDD a_2275_550# 0.07fF
C1072 w_2214_287# VDD 0.22fF
C1073 VDD a_2980_252# 0.07fF
C1074 a_587_n168# a2 0.10fF
C1075 a_1447_n1# a_1252_n84# 0.28fF
C1076 w_2962_470# enb0c 0.06fF
C1077 a_1447_n1# VDD 0.06fF
C1078 VDD enb0c 0.27fF
C1079 gnd b3 0.31fF
C1080 w_3697_n53# pequ 0.07fF
C1081 a1 ena0c 0.01fF
C1082 w_1454_n285# d2 0.10fF
C1083 VDD a_2272_271# 0.07fF
C1084 gnd a_2170_281# 0.35fF
C1085 w_366_n331# a_380_n324# 0.13fF
C1086 a_2107_345# a_2095_345# 0.70fF
C1087 w_366_n130# a_112_n123# 0.07fF
C1088 w_674_n285# a0 0.07fF
C1089 enb3as a_1252_n84# 0.18fF
C1090 a0 a_688_n278# 0.10fF
C1091 enb3as VDD 0.07fF
C1092 ena2a enb2a 0.10fF
C1093 w_1829_n802# enb0a 0.10fF
C1094 a_2210_n2# VDD 0.30fF
C1095 gnd enb3a 0.04fF
C1096 VDD a_2911_n360# 0.06fF
C1097 a_2173_560# VDD 0.07fF
C1098 VDD a_1092_n417# 0.03fF
C1099 a_2098_624# a_2247_620# 0.28fF
C1100 w_3146_n524# x3 0.06fF
C1101 a_2899_n212# a_2882_n234# 0.08fF
C1102 w_2986_n150# x1 0.03fF
C1103 a_1887_n5# a_1252_n84# 1.40fF
C1104 a_1887_n5# VDD 0.28fF
C1105 gnd x0 0.17fF
C1106 gnd w_2967_n625# 0.01fF
C1107 w_2332_303# a_2350_276# 0.09fF
C1108 a_587_n168# a1 0.10fF
C1109 sout2 a_2095_345# 1.20fF
C1110 w_2214_287# a_2207_247# 0.09fF
C1111 w_1713_n424# VDD 0.22fF
C1112 enb3c a_3065_n592# 0.08fF
C1113 a_2898_103# a_2910_103# 0.70fF
C1114 a_1887_n5# w_2115_12# 0.07fF
C1115 w_99_n160# a_112_n178# 0.03fF
C1116 w_2964_n491# VDD 0.10fF
C1117 b0 a_1317_n417# 0.10fF
C1118 ena1c a_2980_252# 0.08fF
C1119 x2 a_3599_n44# 0.08fF
C1120 enb2as a_1748_n4# 0.25fF
C1121 x1 x0 0.87fF
C1122 w_1713_n424# d3 0.10fF
C1123 w_1570_19# enb1as 0.16fF
C1124 gnd enb2a 0.17fF
C1125 a_2210_n2# a_2207_247# 0.51fF
C1126 enb0c ena1c 0.01fF
C1127 gnd a_1748_n4# 0.28fF
C1128 x3 ena3c 0.06fF
C1129 w_3582_n50# x2 0.06fF
C1130 w_2337_858# a_2210_562# 0.03fF
C1131 ena1as d1 0.01fF
C1132 VDD a_831_n145# 0.03fF
C1133 b1 a_1473_n145# 0.10fF
C1134 gnd w_2335_582# 0.23fF
C1135 b3 ena0c 0.01fF
C1136 w_1307_n285# VDD 0.22fF
C1137 enb1c a_2899_n212# 0.08fF
C1138 x3 a_3163_n518# 0.08fF
C1139 w_817_n152# a_831_n145# 0.10fF
C1140 a0 a_693_n145# 0.10fF
C1141 w_2964_n491# a_2977_n509# 0.03fF
C1142 gnd a_380_n354# 0.21fF
C1143 w_3697_n53# VDD 0.25fF
C1144 a_2110_60# ena3as 0.25fF
C1145 a_2244_341# sout2 0.70fF
C1146 a_2173_n4# gnd 0.35fF
C1147 w_2117_852# ena0as 0.09fF
C1148 sout3 a_2210_n2# 0.08fF
C1149 VDD a_3221_530# 0.03fF
C1150 w_670_n424# VDD 0.22fF
C1151 w_1829_n573# and2 0.03fF
C1152 a_2129_19# ena3as 0.04fF
C1153 w_1829_n468# and3 0.03fF
C1154 d2 a2 0.11fF
C1155 VDD a_1326_n145# 0.03fF
C1156 gnd a_3304_n443# 0.03fF
C1157 ena2a enb1a 0.01fF
C1158 ena3a enb0a 0.01fF
C1159 x3 ena2c 0.28fF
C1160 w_2117_852# a_1435_n1# 0.07fF
C1161 a_2098_60# a_2110_60# 0.70fF
C1162 VDD w4 0.07fF
C1163 w_670_n424# d3 0.10fF
C1164 a_587_n168# b3 0.10fF
C1165 VDD ena0a 0.07fF
C1166 a_1584_n3# w_2115_576# 0.07fF
C1167 a_2081_38# ena3as 0.30fF
C1168 w_2985_165# gnd 0.00fF
C1169 w_3473_386# a_2980_319# 0.06fF
C1170 w_2964_n491# ena1c 0.06fF
C1171 gnd a_2210_562# 0.87fF
C1172 a_2218_597# VDD 0.03fF
C1173 VDD a_112_n123# 0.35fF
C1174 w_2223_918# a_2249_896# 0.07fF
C1175 enb0c a_2975_n443# 0.10fF
C1176 w_2221_78# VDD 0.08fF
C1177 gnd ena0as 0.05fF
C1178 gnd a_2883_n80# 0.16fF
C1179 w_3335_424# a_3423_395# 0.02fF
C1180 w_2885_n190# a_2882_n234# 0.12fF
C1181 a_2081_38# a_2098_60# 0.08fF
C1182 b3 enb2c 0.01fF
C1183 VDD x3 0.28fF
C1184 a3 a_1092_n417# 0.10fF
C1185 w_958_n285# ena2c 0.03fF
C1186 w_1459_n152# a_1473_n145# 0.10fF
C1187 a_1435_n1# gnd 0.08fF
C1188 gnd a_2110_624# 0.28fF
C1189 w_1454_n285# b1 0.07fF
C1190 w_3419_n365# VDD 0.32fF
C1191 w_3204_524# x1 0.06fF
C1192 a_3663_329# a_3616_352# 0.02fF
C1193 d2 a1 0.11fF
C1194 ena1a enb1a 0.10fF
C1195 w_1829_n802# ena0a 0.07fF
C1196 gnd a_2078_323# 0.04fF
C1197 gnd enb1a 0.17fF
C1198 w_1722_18# a_1719_n26# 0.12fF
C1199 w_679_n152# a_693_n145# 0.10fF
C1200 w_1194_n68# a_1208_n61# 0.10fF
C1201 gnd b0 0.31fF
C1202 ena2as a_1252_n84# 0.07fF
C1203 ena2as VDD 0.19fF
C1204 w_963_n152# a2 0.07fF
C1205 a_1736_n4# ena3as 0.10fF
C1206 w_2886_n36# a_2883_n80# 0.12fF
C1207 a_1736_n4# a_2095_345# 1.27fF
C1208 w_3654_474# a_3306_495# 0.06fF
C1209 w_2884_125# a_2910_103# 0.07fF
C1210 w_1082_n285# d2 0.10fF
C1211 w_2084_82# a_2110_60# 0.07fF
C1212 x3 a_2977_n509# 0.01fF
C1213 gnd s0 0.26fF
C1214 VDD w_958_n285# 0.22fF
C1215 gnd a_2881_81# 0.16fF
C1216 gnd a_380_n288# 0.28fF
C1217 VDD a_3549_357# 0.09fF
C1218 a_1418_n23# w_1421_21# 0.12fF
C1219 enb0as a_1447_n1# 0.25fF
C1220 w_2885_n190# enb1c 0.16fF
C1221 w_2221_642# sout1 0.13fF
C1222 b3 enb1c 0.01fF
C1223 VDD a_380_n258# 0.11fF
C1224 a2 a_977_n145# 0.10fF
C1225 a_2218_33# a_2210_n2# 0.16fF
C1226 a_2218_597# a_2098_624# 0.14fF
C1227 w_3204_524# ena0c 0.06fF
C1228 gnd a_3436_n359# 0.05fF
C1229 a_2081_38# w_2084_82# 0.12fF
C1230 w_1722_n152# VDD 0.22fF
C1231 gnd a_1317_n417# 0.03fF
C1232 x3 ena1c 0.24fF
C1233 d2 a_3711_n46# 0.24fF
C1234 VDD a_2911_n212# 0.06fF
C1235 sout3 w_2221_78# 0.13fF
C1236 a_2275_550# w_2217_566# 0.03fF
C1237 a2 a_972_n278# 0.10fF
C1238 gnd a_1612_n145# 0.03fF
C1239 w_2332_303# a_2272_271# 0.11fF
C1240 a_2083_878# ena0as 0.30fF
C1241 d2 b3 0.11fF
C1242 x1 a_3436_n359# 0.08fF
C1243 w_2086_922# a_2112_900# 0.07fF
C1244 w_1312_n152# b0 0.07fF
C1245 gnd a_3490_392# 0.03fF
C1246 a_2129_583# VDD 0.03fF
C1247 b0 ena0c 0.01fF
C1248 w_3645_n306# w4 0.06fF
C1249 w_2332_303# a_2210_n2# 0.03fF
C1250 w_1194_n68# a_1252_n84# 0.03fF
C1251 VDD a_2977_386# 0.08fF
C1252 w_1194_n68# VDD 0.22fF
C1253 a_1435_n1# a_2083_878# 0.14fF
C1254 w_1082_n285# a_1096_n278# 0.10fF
C1255 ena0as a_587_n168# 0.01fF
C1256 a_2228_294# VDD 0.03fF
C1257 and0 Gnd 0.06fF
C1258 a_1843_n795# Gnd 0.33fF
C1259 and1 Gnd 0.06fF
C1260 a_1843_n688# Gnd 0.33fF
C1261 a_3065_n592# Gnd 0.36fF
C1262 a_2980_n643# Gnd 0.81fF
C1263 a_3163_n518# Gnd 0.41fF
C1264 a_2980_n576# Gnd 1.68fF
C1265 a_3304_n443# Gnd 0.44fF
C1266 a_2977_n509# Gnd 2.41fF
C1267 a_3436_n359# Gnd 0.51fF
C1268 a_2975_n443# Gnd 3.44fF
C1269 a_2911_n360# Gnd 0.27fF
C1270 lsr Gnd 0.08fF
C1271 a_3661_n330# Gnd 0.35fF
C1272 w4 Gnd 6.09fF
C1273 w3 Gnd 1.09fF
C1274 w2 Gnd 3.09fF
C1275 w1 Gnd 1.42fF
C1276 a_2882_n382# Gnd 1.87fF
C1277 a_2899_n360# Gnd 1.11fF
C1278 a_2911_n212# Gnd 0.27fF
C1279 a_2882_n234# Gnd 1.87fF
C1280 a_2899_n212# Gnd 1.11fF
C1281 equ Gnd 0.06fF
C1282 a_3711_n46# Gnd 0.40fF
C1283 pequ Gnd 0.31fF
C1284 a_3599_n44# Gnd 0.44fF
C1285 x0 Gnd 3.41fF
C1286 a_3616_352# Gnd 0.36fF
C1287 a_2912_n58# Gnd 0.27fF
C1288 a_2883_n80# Gnd 1.87fF
C1289 a_2900_n58# Gnd 1.11fF
C1290 a_2910_103# Gnd 0.27fF
C1291 a_2881_81# Gnd 1.87fF
C1292 a_2898_103# Gnd 1.11fF
C1293 a_2980_252# Gnd 3.37fF
C1294 a_3490_392# Gnd 0.41fF
C1295 a_2980_319# Gnd 1.99fF
C1296 gtr Gnd 0.08fF
C1297 a_3670_450# Gnd 0.35fF
C1298 a_3663_329# Gnd 1.10fF
C1299 a_3549_357# Gnd 1.65fF
C1300 a_3423_395# Gnd 2.26fF
C1301 a_3352_430# Gnd 0.44fF
C1302 a_2977_386# Gnd 3.09fF
C1303 and2 Gnd 0.06fF
C1304 a_1843_n566# Gnd 0.33fF
C1305 and3 Gnd 0.06fF
C1306 a_1843_n461# Gnd 0.33fF
C1307 enb3a Gnd 0.86fF
C1308 a_1727_n417# Gnd 0.33fF
C1309 enb2a Gnd 2.12fF
C1310 a_1603_n417# Gnd 0.33fF
C1311 enb1a Gnd 3.65fF
C1312 a_1464_n417# Gnd 0.33fF
C1313 enb0a Gnd 5.12fF
C1314 a_1317_n417# Gnd 0.33fF
C1315 ena3a Gnd 8.53fF
C1316 a_1092_n417# Gnd 0.33fF
C1317 ena2a Gnd 11.09fF
C1318 a_968_n417# Gnd 0.33fF
C1319 ena1a Gnd 14.13fF
C1320 a_822_n417# Gnd 0.33fF
C1321 ena0a Gnd 9.02fF
C1322 a_684_n417# Gnd 0.33fF
C1323 enb3c Gnd 9.55fF
C1324 a_1731_n278# Gnd 0.33fF
C1325 enb2c Gnd 14.17fF
C1326 a_1607_n278# Gnd 0.33fF
C1327 enb1c Gnd 16.69fF
C1328 a_1468_n278# Gnd 0.33fF
C1329 a_1321_n278# Gnd 0.33fF
C1330 ena3c Gnd 26.03fF
C1331 a_1096_n278# Gnd 0.33fF
C1332 ena2c Gnd 26.33fF
C1333 a_972_n278# Gnd 0.33fF
C1334 a_380_n354# Gnd 0.10fF
C1335 d3 Gnd 11.15fF
C1336 a_380_n324# Gnd 0.40fF
C1337 ena1c Gnd 25.57fF
C1338 a_826_n278# Gnd 0.33fF
C1339 a_380_n288# Gnd 0.10fF
C1340 a_688_n278# Gnd 0.33fF
C1341 enb0c Gnd 18.65fF
C1342 a_3306_495# Gnd 3.38fF
C1343 a_3221_530# Gnd 0.51fF
C1344 x1 Gnd 13.78fF
C1345 x2 Gnd 16.95fF
C1346 x3 Gnd 22.96fF
C1347 ena0c Gnd 29.31fF
C1348 a_2975_452# Gnd 2.16fF
C1349 a_380_n258# Gnd 0.40fF
C1350 a_380_n222# Gnd 0.10fF
C1351 a_380_n192# Gnd 0.40fF
C1352 a_1736_n145# Gnd 0.33fF
C1353 b3 Gnd 4.34fF
C1354 a_1612_n145# Gnd 0.33fF
C1355 b2 Gnd 4.53fF
C1356 a_1473_n145# Gnd 0.33fF
C1357 b1 Gnd 4.52fF
C1358 a_1326_n145# Gnd 0.33fF
C1359 b0 Gnd 4.65fF
C1360 a_1101_n145# Gnd 0.33fF
C1361 a3 Gnd 4.48fF
C1362 a_977_n145# Gnd 0.33fF
C1363 a2 Gnd 4.57fF
C1364 a_831_n145# Gnd 0.33fF
C1365 a1 Gnd 4.60fF
C1366 a_693_n145# Gnd 0.33fF
C1367 a0 Gnd 4.71fF
C1368 a_547_n182# Gnd 0.31fF
C1369 a_380_n153# Gnd 0.10fF
C1370 s1 Gnd 2.33fF
C1371 d0 Gnd 1.36fF
C1372 a_380_n123# Gnd 0.40fF
C1373 a_112_n178# Gnd 2.70fF
C1374 a_112_n123# Gnd 4.39fF
C1375 s0 Gnd 5.75fF
C1376 a_1208_n61# Gnd 0.33fF
C1377 a_587_n168# Gnd 10.28fF
C1378 d1 Gnd 6.26fF
C1379 a_2231_9# Gnd 0.33fF
C1380 cout Gnd 0.12fF
C1381 a_2129_19# Gnd 0.33fF
C1382 a_1899_n5# Gnd 0.27fF
C1383 a_2353_n9# Gnd 0.31fF
C1384 a_2173_n4# Gnd 2.37fF
C1385 a_2275_n14# Gnd 1.10fF
C1386 a_2247_56# Gnd 0.27fF
C1387 sout3 Gnd 0.24fF
C1388 a_2110_60# Gnd 0.27fF
C1389 a_2098_60# Gnd 3.48fF
C1390 a_1887_n5# Gnd 3.22fF
C1391 a_2218_33# Gnd 1.88fF
C1392 ena3as Gnd 3.02fF
C1393 enb3as Gnd 3.33fF
C1394 a_1748_n4# Gnd 0.27fF
C1395 a_1870_n27# Gnd 1.87fF
C1396 enb2as Gnd 2.94fF
C1397 a_1596_n3# Gnd 0.27fF
C1398 a_1719_n26# Gnd 1.87fF
C1399 enb1as Gnd 2.87fF
C1400 a_1447_n1# Gnd 0.27fF
C1401 a_1567_n25# Gnd 1.87fF
C1402 enb0as Gnd 2.90fF
C1403 a_1418_n23# Gnd 1.87fF
C1404 a_2081_38# Gnd 1.87fF
C1405 a_2228_294# Gnd 0.33fF
C1406 a_2210_n2# Gnd 5.24fF
C1407 a_2126_304# Gnd 0.33fF
C1408 a_2350_276# Gnd 0.31fF
C1409 a_2170_281# Gnd 2.37fF
C1410 a_2272_271# Gnd 1.10fF
C1411 a_2244_341# Gnd 0.27fF
C1412 sout2 Gnd 0.24fF
C1413 a_2107_345# Gnd 0.27fF
C1414 a_2095_345# Gnd 3.48fF
C1415 a_1736_n4# Gnd 7.71fF
C1416 a_2215_318# Gnd 1.88fF
C1417 ena2as Gnd 3.04fF
C1418 a_2078_323# Gnd 1.87fF
C1419 d2 Gnd 31.97fF
C1420 a_2231_573# Gnd 0.33fF
C1421 a_2207_247# Gnd 4.21fF
C1422 a_2129_583# Gnd 0.33fF
C1423 a_2353_555# Gnd 0.31fF
C1424 a_2173_560# Gnd 2.37fF
C1425 a_2275_550# Gnd 1.10fF
C1426 a_2247_620# Gnd 0.27fF
C1427 sout1 Gnd 0.24fF
C1428 a_2110_624# Gnd 0.27fF
C1429 a_2098_624# Gnd 3.48fF
C1430 a_1584_n3# Gnd 12.41fF
C1431 a_2218_597# Gnd 1.88fF
C1432 ena1as Gnd 3.46fF
C1433 a_2081_602# Gnd 1.87fF
C1434 a_2233_849# Gnd 0.33fF
C1435 a_2210_562# Gnd 5.92fF
C1436 a_2131_859# Gnd 0.33fF
C1437 a_2355_831# Gnd 0.31fF
C1438 a_2175_836# Gnd 2.37fF
C1439 a_2277_826# Gnd 1.10fF
C1440 a_2249_896# Gnd 0.27fF
C1441 sout0 Gnd 0.24fF
C1442 a_1252_n84# Gnd 11.54fF
C1443 gnd Gnd 63.97fF
C1444 VDD Gnd 82.24fF
C1445 a_2112_900# Gnd 0.27fF
C1446 a_2100_900# Gnd 3.48fF
C1447 a_1435_n1# Gnd 17.15fF
C1448 a_2220_873# Gnd 1.88fF
C1449 ena0as Gnd 4.63fF
C1450 a_2083_878# Gnd 1.87fF
C1451 w_1829_n802# Gnd 1.48fF
C1452 w_1829_n695# Gnd 1.48fF
C1453 w_2967_n625# Gnd 0.48fF
C1454 w_3051_n599# Gnd 1.54fF
C1455 w_2967_n558# Gnd 0.48fF
C1456 w_1829_n573# Gnd 1.48fF
C1457 w_3146_n524# Gnd 2.10fF
C1458 w_2964_n491# Gnd 0.48fF
C1459 w_3287_n449# Gnd 2.38fF
C1460 w_1829_n468# Gnd 1.48fF
C1461 w_2962_n425# Gnd 0.48fF
C1462 w_1713_n424# Gnd 1.48fF
C1463 w_1589_n424# Gnd 1.48fF
C1464 w_1450_n424# Gnd 1.48fF
C1465 w_1303_n424# Gnd 1.48fF
C1466 w_1078_n424# Gnd 1.48fF
C1467 w_954_n424# Gnd 1.48fF
C1468 w_808_n424# Gnd 1.48fF
C1469 w_670_n424# Gnd 1.48fF
C1470 w_3419_n365# Gnd 2.70fF
C1471 w_2885_n338# Gnd 2.10fF
C1472 w_366_n331# Gnd 1.62fF
C1473 w_3645_n306# Gnd 1.88fF
C1474 w_2986_n298# Gnd 0.48fF
C1475 w_1717_n285# Gnd 1.48fF
C1476 w_1593_n285# Gnd 1.48fF
C1477 w_1454_n285# Gnd 1.48fF
C1478 w_1307_n285# Gnd 1.48fF
C1479 w_1082_n285# Gnd 1.48fF
C1480 w_958_n285# Gnd 1.48fF
C1481 w_812_n285# Gnd 1.48fF
C1482 w_674_n285# Gnd 1.48fF
C1483 w_366_n265# Gnd 1.62fF
C1484 w_2885_n190# Gnd 2.10fF
C1485 w_366_n199# Gnd 1.61fF
C1486 w_2986_n150# Gnd 0.48fF
C1487 w_1722_n152# Gnd 1.48fF
C1488 w_1598_n152# Gnd 1.48fF
C1489 w_1459_n152# Gnd 1.48fF
C1490 w_1312_n152# Gnd 1.48fF
C1491 w_1087_n152# Gnd 1.48fF
C1492 w_963_n152# Gnd 1.48fF
C1493 w_817_n152# Gnd 1.48fF
C1494 w_679_n152# Gnd 1.48fF
C1495 w_529_n155# Gnd 1.56fF
C1496 w_99_n160# Gnd 0.48fF
C1497 w_366_n130# Gnd 1.62fF
C1498 w_99_n105# Gnd 0.48fF
C1499 w_3697_n53# Gnd 1.77fF
C1500 w_3582_n50# Gnd 2.38fF
C1501 w_1194_n68# Gnd 1.48fF
C1502 w_2886_n36# Gnd 2.10fF
C1503 w_2987_4# Gnd 0.48fF
C1504 w_2217_2# Gnd 1.48fF
C1505 w_2335_18# Gnd 1.56fF
C1506 w_2115_12# Gnd 1.48fF
C1507 w_1873_17# Gnd 2.10fF
C1508 w_1722_18# Gnd 2.10fF
C1509 w_1570_19# Gnd 2.10fF
C1510 w_1421_21# Gnd 2.10fF
C1511 w_2221_78# Gnd 2.10fF
C1512 w_2084_82# Gnd 2.10fF
C1513 w_2884_125# Gnd 2.10fF
C1514 w_2985_165# Gnd 0.48fF
C1515 w_2967_270# Gnd 0.48fF
C1516 w_2214_287# Gnd 1.48fF
C1517 w_2332_303# Gnd 1.56fF
C1518 w_2112_297# Gnd 1.48fF
C1519 w_3602_345# Gnd 1.54fF
C1520 w_2967_337# Gnd 0.48fF
C1521 w_2218_363# Gnd 2.10fF
C1522 w_3473_386# Gnd 2.10fF
C1523 w_2081_367# Gnd 2.10fF
C1524 w_2964_404# Gnd 0.48fF
C1525 w_3335_424# Gnd 2.38fF
C1526 w_3654_474# Gnd 1.88fF
C1527 w_2962_470# Gnd 0.48fF
C1528 w_3204_524# Gnd 2.70fF
C1529 w_2217_566# Gnd 1.48fF
C1530 w_2335_582# Gnd 1.56fF
C1531 w_2115_576# Gnd 1.48fF
C1532 w_2221_642# Gnd 2.10fF
C1533 w_2084_646# Gnd 2.10fF
C1534 w_2219_842# Gnd 1.48fF
C1535 w_2337_858# Gnd 1.56fF
C1536 w_2117_852# Gnd 1.48fF
C1537 w_2223_918# Gnd 2.10fF
C1538 w_2086_922# Gnd 2.10fF


* Vi1 s0 gnd pulse(1.8 0 10n 100p 100p 200n 400n)
* Vi2 s1 gnd pulse(1.8 0 10n 100p 100p 200n 400n)
* Vi1 s0 gnd pulse(0 1.8 10n 100p 100p 200n 400n)
* Vi2 s1 gnd pulse(0 1.8 10n 100p 100p 200n 400n)

* Vi1 s0 gnd DC SUPPLY
Vi2 s1 gnd DC 0
Vi1 s0 gnd DC 0
* Vi2 s1 gnd DC 0



* V_a0 a0 gnd pulse(0 1.8 0ns 100ps 799ns 800ns)
* V_a0 a0 gnd pulse(1.8 0 0ns 100ps 799ns 800ns)
* V_a1 a1 gnd pulse(1.8 0 0ns 100ps 799ns 800ns)
* V_a1 a1 gnd pulse(0 1.8 0ns 100ps 799ns 800ns)
* V_a2 a2 gnd pulse(0 1.8 0ns 100ps 799ns 800ns)
* V_a2 a2 gnd pulse(1.8 0 0ns 100ps 799ns 800ns)
* V_a3 a3 gnd pulse(0 1.8 0ns 100ps 799ns 800ns)
* V_a3 a3 gnd pulse(1.8 0 0ns 100ps 799ns 800ns)
* V_b0 b0 gnd pulse(0 1.8 0ns 100ps 799ns 800ns)
* V_b0 b0 gnd pulse(1.8 0 0ns 100ps 799ns 800ns)
* V_b1 b1 gnd pulse(1.8 0 0ns 100ps 799ns 800ns)
* V_b1 b1 gnd pulse(0 1.8 0ns 100ps 799ns 800ns)
* V_b2 b2 gnd pulse(0 1.8 0ns 100ps 799ns 800ns)
* V_b2 b2 gnd pulse(1.8 0 0ns 100ps 799ns 800ns)
* V_b3 b3 gnd pulse(0 1.8 0ns 100ps 799ns 800ns)
* V_b3 b3 gnd pulse(1.8 0 0ns 100ps 799ns 800ns)


* V_a0 a0 gnd PULSE(0 1.8 0ns 100ps 100ps 100ns 400ns)
* V_a1 a1 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 600ns)
* V_a2 a2 gnd PULSE(0 1.8 0ns 100ps 100ps 400ns 800ns)
* V_a3 a3 gnd PULSE(0 1.8 0ns 100ps 100ps 200ns 400ns)
* V_b0 b0 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 600ns)
* V_b1 b1 gnd PULSE(0 1.8 0ns 100ps 100ps 100ns 800ns)
* V_b2 b2 gnd PULSE(0 1.8 0ns 100ps 100ps 200ns 400ns)
* V_b3 b3 gnd PULSE(0 1.8 0ns 100ps 100ps 400ns 800ns)

V_b0 b0 gnd pulse(0 1.8 0n 100p 100p 200n 400n)
V_b1 b1 gnd pulse(0 1.8 0n 100p 100p 200n 400n)
V_b2 b2 gnd pulse(0 1.8 0n 100p 100p 200n 400n)
V_b3 b3 gnd pulse(0 1.8 0n 100p 100p 200n 400n)
V_a0 a0 gnd DC 0
V_a1 a1 gnd DC 0
V_a2 a2 gnd DC 0
V_a3 a3 gnd DC 0

V1 VDD gnd 1.8


.tran 1n 810n

*target text

.control
run
* set color0 = rgb:f/f/e
* set color1 = black
* plot v(s0) v(s1)+2 v(d0)+4 v(d1)+6 v(d2)+8 v(d3)+10 title "Select lines"
* plot v(a0) v(a1)+2 v(a2)+4 v(a3)+6 v(b0)+8 v(b1)+10 v(b2)+12 v(b3)+14 title "inputs"
* plot v(ena0as) v(ena1as)+2 v(ena2as)+4 v(ena3as)+6 v(enb0as)+8 v(enb1as)+10 v(enb2as)+12 v(enb3as)+14 title "adder enable"
* plot v(ena0c) v(ena1c)+2 v(ena2c)+4 v(ena3c)+6 v(enb0c)+8 v(enb1c)+10 v(enb2c)+12 v(enb3c)+14 title "comp enable"
* plot v(ena0a) v(ena1a)+2 v(ena2a)+4 v(ena3a)+6 v(enb0a)+8 v(enb1a)+10 v(enb2a)+12 v(enb3a)+14 title "and enable"
* plot v(and0) v(and1)+2 v(and2)+4 v(and3)+6 title "ander"
* plot v(gtr) v(equ)+2 v(lsr)+4 title "comaparator"
* plot v(sout0) v(sout1)+2 v(sout2)+4 v(sout3)+6 v(cout)+8 title "adder/ subtractor"
quit
.end
.endc