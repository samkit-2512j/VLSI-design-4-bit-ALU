magic
tech scmos
timestamp 1701518043
<< nwell >>
rect 2086 922 2177 945
rect 2223 918 2314 941
rect 2117 852 2187 873
rect 2337 863 2407 882
rect 2219 842 2289 863
rect 2337 858 2382 863
rect 2084 646 2175 669
rect 2221 642 2312 665
rect 2115 576 2185 597
rect 2335 587 2405 606
rect 2217 566 2287 587
rect 2335 582 2380 587
rect 3204 524 3321 547
rect 2962 470 2987 489
rect 3654 474 3743 495
rect 3335 424 3438 447
rect 2964 404 2989 423
rect 2081 367 2172 390
rect 3473 386 3564 409
rect 2218 363 2309 386
rect 2967 337 2992 356
rect 3602 345 3675 366
rect 2112 297 2182 318
rect 2332 308 2402 327
rect 2214 287 2284 308
rect 2332 303 2377 308
rect 2967 270 2992 289
rect 2985 165 3010 184
rect 2884 125 2975 148
rect 2084 82 2175 105
rect 2221 78 2312 101
rect 1421 21 1512 44
rect 1570 19 1661 42
rect 1722 18 1813 41
rect 1873 17 1964 40
rect 2115 12 2185 33
rect 2335 23 2405 42
rect 2217 2 2287 23
rect 2335 18 2380 23
rect 2987 4 3012 23
rect 2886 -36 2977 -13
rect 1194 -68 1264 -47
rect 3582 -50 3685 -27
rect 3697 -53 3781 -32
rect 99 -105 124 -86
rect 366 -128 445 -109
rect 366 -130 420 -128
rect 99 -160 124 -141
rect 529 -150 599 -131
rect 529 -155 574 -150
rect 679 -152 749 -131
rect 817 -152 887 -131
rect 963 -152 1033 -131
rect 1087 -152 1157 -131
rect 1312 -152 1382 -131
rect 1459 -152 1529 -131
rect 1598 -152 1668 -131
rect 1722 -152 1792 -131
rect 2986 -150 3011 -131
rect 368 -181 445 -178
rect 366 -197 445 -181
rect 2885 -190 2976 -167
rect 366 -199 420 -197
rect 366 -263 445 -244
rect 366 -265 420 -263
rect 674 -285 744 -264
rect 812 -285 882 -264
rect 958 -285 1028 -264
rect 1082 -285 1152 -264
rect 1307 -285 1377 -264
rect 1454 -285 1524 -264
rect 1593 -285 1663 -264
rect 1717 -285 1787 -264
rect 2986 -298 3011 -279
rect 3645 -306 3734 -285
rect 366 -329 445 -310
rect 366 -331 420 -329
rect 2885 -338 2976 -315
rect 3419 -365 3536 -342
rect 670 -424 740 -403
rect 808 -424 878 -403
rect 954 -424 1024 -403
rect 1078 -424 1148 -403
rect 1303 -424 1373 -403
rect 1450 -424 1520 -403
rect 1589 -424 1659 -403
rect 1713 -424 1783 -403
rect 2962 -425 2987 -406
rect 1829 -468 1899 -447
rect 3287 -449 3390 -426
rect 2964 -491 2989 -472
rect 3146 -524 3237 -501
rect 1829 -573 1899 -552
rect 2967 -558 2992 -539
rect 3051 -599 3124 -578
rect 2967 -625 2992 -606
rect 1829 -695 1899 -674
rect 1829 -802 1899 -781
<< ntransistor >>
rect 2098 900 2100 905
rect 2117 900 2119 905
rect 2142 900 2144 905
rect 2161 900 2163 905
rect 2235 896 2237 901
rect 2254 896 2256 901
rect 2279 896 2281 901
rect 2298 896 2300 901
rect 2173 836 2175 840
rect 2129 829 2131 836
rect 2144 829 2146 836
rect 2393 845 2395 849
rect 2353 831 2355 840
rect 2362 831 2364 840
rect 2275 826 2277 830
rect 2231 819 2233 826
rect 2246 819 2248 826
rect 2096 624 2098 629
rect 2115 624 2117 629
rect 2140 624 2142 629
rect 2159 624 2161 629
rect 2233 620 2235 625
rect 2252 620 2254 625
rect 2277 620 2279 625
rect 2296 620 2298 625
rect 2171 560 2173 564
rect 2127 553 2129 560
rect 2142 553 2144 560
rect 2391 569 2393 573
rect 2351 555 2353 564
rect 2360 555 2362 564
rect 2273 550 2275 554
rect 2229 543 2231 550
rect 2244 543 2246 550
rect 2093 345 2095 350
rect 2112 345 2114 350
rect 2137 345 2139 350
rect 2156 345 2158 350
rect 2230 341 2232 346
rect 2249 341 2251 346
rect 2274 341 2276 346
rect 2293 341 2295 346
rect 2168 281 2170 285
rect 2124 274 2126 281
rect 2139 274 2141 281
rect 2388 290 2390 294
rect 2348 276 2350 285
rect 2357 276 2359 285
rect 2270 271 2272 275
rect 2226 264 2228 271
rect 2241 264 2243 271
rect 1433 -1 1435 4
rect 1452 -1 1454 4
rect 1477 -1 1479 4
rect 1496 -1 1498 4
rect 1582 -3 1584 2
rect 1601 -3 1603 2
rect 1626 -3 1628 2
rect 1645 -3 1647 2
rect 1734 -4 1736 1
rect 1753 -4 1755 1
rect 1778 -4 1780 1
rect 1797 -4 1799 1
rect 2096 60 2098 65
rect 2115 60 2117 65
rect 2140 60 2142 65
rect 2159 60 2161 65
rect 2233 56 2235 61
rect 2252 56 2254 61
rect 2277 56 2279 61
rect 2296 56 2298 61
rect 1885 -5 1887 0
rect 1904 -5 1906 0
rect 1929 -5 1931 0
rect 1948 -5 1950 0
rect 2171 -4 2173 0
rect 2127 -11 2129 -4
rect 2142 -11 2144 -4
rect 2391 5 2393 9
rect 2351 -9 2353 0
rect 2360 -9 2362 0
rect 2273 -14 2275 -10
rect 2229 -21 2231 -14
rect 2244 -21 2246 -14
rect 110 -123 112 -119
rect 431 -146 433 -142
rect 378 -153 380 -146
rect 404 -153 406 -146
rect 1250 -84 1252 -80
rect 1206 -91 1208 -84
rect 1221 -91 1223 -84
rect 585 -168 587 -164
rect 735 -168 737 -164
rect 873 -168 875 -164
rect 1019 -168 1021 -164
rect 1143 -168 1145 -164
rect 1368 -168 1370 -164
rect 1515 -168 1517 -164
rect 1654 -168 1656 -164
rect 1778 -168 1780 -164
rect 110 -178 112 -174
rect 545 -182 547 -173
rect 554 -182 556 -173
rect 691 -175 693 -168
rect 706 -175 708 -168
rect 829 -175 831 -168
rect 844 -175 846 -168
rect 975 -175 977 -168
rect 990 -175 992 -168
rect 1099 -175 1101 -168
rect 1114 -175 1116 -168
rect 1324 -175 1326 -168
rect 1339 -175 1341 -168
rect 1471 -175 1473 -168
rect 1486 -175 1488 -168
rect 1610 -175 1612 -168
rect 1625 -175 1627 -168
rect 1734 -175 1736 -168
rect 1749 -175 1751 -168
rect 431 -215 433 -211
rect 378 -222 380 -215
rect 404 -222 406 -215
rect 3219 495 3221 505
rect 3234 495 3236 505
rect 3249 495 3251 505
rect 3264 495 3266 505
rect 3278 495 3280 505
rect 3304 495 3306 505
rect 431 -281 433 -277
rect 378 -288 380 -281
rect 404 -288 406 -281
rect 730 -301 732 -297
rect 686 -308 688 -301
rect 701 -308 703 -301
rect 431 -347 433 -343
rect 378 -354 380 -347
rect 404 -354 406 -347
rect 868 -301 870 -297
rect 824 -308 826 -301
rect 839 -308 841 -301
rect 1014 -301 1016 -297
rect 970 -308 972 -301
rect 985 -308 987 -301
rect 1138 -301 1140 -297
rect 1094 -308 1096 -301
rect 1109 -308 1111 -301
rect 1363 -301 1365 -297
rect 1319 -308 1321 -301
rect 1334 -308 1336 -301
rect 1510 -301 1512 -297
rect 1466 -308 1468 -301
rect 1481 -308 1483 -301
rect 1649 -301 1651 -297
rect 1605 -308 1607 -301
rect 1620 -308 1622 -301
rect 1773 -301 1775 -297
rect 1729 -308 1731 -301
rect 1744 -308 1746 -301
rect 726 -440 728 -436
rect 682 -447 684 -440
rect 697 -447 699 -440
rect 864 -440 866 -436
rect 1010 -440 1012 -436
rect 1134 -440 1136 -436
rect 1359 -440 1361 -436
rect 820 -447 822 -440
rect 835 -447 837 -440
rect 966 -447 968 -440
rect 981 -447 983 -440
rect 1090 -447 1092 -440
rect 1105 -447 1107 -440
rect 1315 -447 1317 -440
rect 1330 -447 1332 -440
rect 1506 -440 1508 -436
rect 1462 -447 1464 -440
rect 1477 -447 1479 -440
rect 1645 -440 1647 -436
rect 1601 -447 1603 -440
rect 1616 -447 1618 -440
rect 1769 -440 1771 -436
rect 1725 -447 1727 -440
rect 1740 -447 1742 -440
rect 1885 -484 1887 -480
rect 1841 -491 1843 -484
rect 1856 -491 1858 -484
rect 2973 452 2975 456
rect 3668 450 3670 457
rect 3680 450 3682 457
rect 3695 450 3697 457
rect 3705 450 3707 457
rect 3728 450 3730 457
rect 3350 395 3352 405
rect 3365 395 3367 405
rect 3385 395 3387 405
rect 3395 395 3397 405
rect 3421 395 3423 405
rect 2975 386 2977 390
rect 2978 319 2980 323
rect 2978 252 2980 256
rect 2996 147 2998 151
rect 2896 103 2898 108
rect 2915 103 2917 108
rect 2940 103 2942 108
rect 2959 103 2961 108
rect 2998 -14 3000 -10
rect 2898 -58 2900 -53
rect 2917 -58 2919 -53
rect 2942 -58 2944 -53
rect 2961 -58 2963 -53
rect 3488 357 3490 367
rect 3503 357 3505 367
rect 3523 357 3525 367
rect 3547 357 3549 367
rect 3661 329 3663 333
rect 3614 322 3616 329
rect 3635 322 3637 329
rect 3767 -69 3769 -65
rect 3597 -79 3599 -69
rect 3612 -79 3614 -69
rect 3632 -79 3634 -69
rect 3642 -79 3644 -69
rect 3668 -79 3670 -69
rect 3709 -76 3711 -69
rect 3735 -76 3737 -69
rect 2997 -168 2999 -164
rect 2897 -212 2899 -207
rect 2916 -212 2918 -207
rect 2941 -212 2943 -207
rect 2960 -212 2962 -207
rect 2997 -316 2999 -312
rect 3659 -330 3661 -323
rect 3671 -330 3673 -323
rect 3686 -330 3688 -323
rect 3696 -330 3698 -323
rect 3719 -330 3721 -323
rect 2897 -360 2899 -355
rect 2916 -360 2918 -355
rect 2941 -360 2943 -355
rect 2960 -360 2962 -355
rect 3434 -394 3436 -384
rect 3449 -394 3451 -384
rect 3464 -394 3466 -384
rect 3479 -394 3481 -384
rect 3493 -394 3495 -384
rect 3519 -394 3521 -384
rect 2973 -443 2975 -439
rect 3302 -478 3304 -468
rect 3317 -478 3319 -468
rect 3337 -478 3339 -468
rect 3347 -478 3349 -468
rect 3373 -478 3375 -468
rect 2975 -509 2977 -505
rect 3161 -553 3163 -543
rect 3176 -553 3178 -543
rect 3196 -553 3198 -543
rect 3220 -553 3222 -543
rect 2978 -576 2980 -572
rect 1885 -589 1887 -585
rect 1841 -596 1843 -589
rect 1856 -596 1858 -589
rect 3110 -615 3112 -611
rect 3063 -622 3065 -615
rect 3084 -622 3086 -615
rect 2978 -643 2980 -639
rect 1885 -711 1887 -707
rect 1841 -718 1843 -711
rect 1856 -718 1858 -711
rect 1885 -818 1887 -814
rect 1841 -825 1843 -818
rect 1856 -825 1858 -818
<< ptransistor >>
rect 2098 931 2100 936
rect 2117 931 2119 936
rect 2142 931 2144 936
rect 2161 931 2163 936
rect 2235 927 2237 932
rect 2254 927 2256 932
rect 2279 927 2281 932
rect 2298 927 2300 932
rect 2353 864 2355 873
rect 2362 864 2364 873
rect 2393 869 2395 873
rect 2129 859 2131 864
rect 2144 859 2146 864
rect 2173 860 2175 864
rect 2231 849 2233 854
rect 2246 849 2248 854
rect 2275 850 2277 854
rect 2096 655 2098 660
rect 2115 655 2117 660
rect 2140 655 2142 660
rect 2159 655 2161 660
rect 2233 651 2235 656
rect 2252 651 2254 656
rect 2277 651 2279 656
rect 2296 651 2298 656
rect 2351 588 2353 597
rect 2360 588 2362 597
rect 2391 593 2393 597
rect 2127 583 2129 588
rect 2142 583 2144 588
rect 2171 584 2173 588
rect 2229 573 2231 578
rect 2244 573 2246 578
rect 2273 574 2275 578
rect 2093 376 2095 381
rect 2112 376 2114 381
rect 2137 376 2139 381
rect 2156 376 2158 381
rect 2230 372 2232 377
rect 2249 372 2251 377
rect 2274 372 2276 377
rect 2293 372 2295 377
rect 2348 309 2350 318
rect 2357 309 2359 318
rect 2388 314 2390 318
rect 2124 304 2126 309
rect 2139 304 2141 309
rect 2168 305 2170 309
rect 2226 294 2228 299
rect 2241 294 2243 299
rect 2270 295 2272 299
rect 1433 30 1435 35
rect 1452 30 1454 35
rect 1477 30 1479 35
rect 1496 30 1498 35
rect 1582 28 1584 33
rect 1601 28 1603 33
rect 1626 28 1628 33
rect 1645 28 1647 33
rect 1734 27 1736 32
rect 1753 27 1755 32
rect 1778 27 1780 32
rect 1797 27 1799 32
rect 2096 91 2098 96
rect 2115 91 2117 96
rect 2140 91 2142 96
rect 2159 91 2161 96
rect 2233 87 2235 92
rect 2252 87 2254 92
rect 2277 87 2279 92
rect 2296 87 2298 92
rect 1885 26 1887 31
rect 1904 26 1906 31
rect 1929 26 1931 31
rect 1948 26 1950 31
rect 2351 24 2353 33
rect 2360 24 2362 33
rect 2391 29 2393 33
rect 2127 19 2129 24
rect 2142 19 2144 24
rect 2171 20 2173 24
rect 2229 9 2231 14
rect 2244 9 2246 14
rect 2273 10 2275 14
rect 1206 -61 1208 -56
rect 1221 -61 1223 -56
rect 1250 -60 1252 -56
rect 110 -99 112 -95
rect 378 -123 380 -118
rect 404 -123 406 -118
rect 431 -122 433 -118
rect 110 -154 112 -150
rect 545 -149 547 -140
rect 554 -149 556 -140
rect 585 -144 587 -140
rect 691 -145 693 -140
rect 706 -145 708 -140
rect 735 -144 737 -140
rect 829 -145 831 -140
rect 844 -145 846 -140
rect 873 -144 875 -140
rect 975 -145 977 -140
rect 990 -145 992 -140
rect 1019 -144 1021 -140
rect 1099 -145 1101 -140
rect 1114 -145 1116 -140
rect 1143 -144 1145 -140
rect 1324 -145 1326 -140
rect 1339 -145 1341 -140
rect 1368 -144 1370 -140
rect 1471 -145 1473 -140
rect 1486 -145 1488 -140
rect 1515 -144 1517 -140
rect 1610 -145 1612 -140
rect 1625 -145 1627 -140
rect 1654 -144 1656 -140
rect 1734 -145 1736 -140
rect 1749 -145 1751 -140
rect 1778 -144 1780 -140
rect 378 -192 380 -187
rect 404 -192 406 -187
rect 431 -191 433 -187
rect 378 -258 380 -253
rect 404 -258 406 -253
rect 431 -257 433 -253
rect 3219 530 3221 540
rect 3234 530 3236 540
rect 3249 530 3251 540
rect 3264 530 3266 540
rect 3278 530 3280 540
rect 3304 530 3306 540
rect 2973 476 2975 480
rect 686 -278 688 -273
rect 701 -278 703 -273
rect 730 -277 732 -273
rect 824 -278 826 -273
rect 839 -278 841 -273
rect 868 -277 870 -273
rect 378 -324 380 -319
rect 404 -324 406 -319
rect 431 -323 433 -319
rect 970 -278 972 -273
rect 985 -278 987 -273
rect 1014 -277 1016 -273
rect 1094 -278 1096 -273
rect 1109 -278 1111 -273
rect 1138 -277 1140 -273
rect 1319 -278 1321 -273
rect 1334 -278 1336 -273
rect 1363 -277 1365 -273
rect 1466 -278 1468 -273
rect 1481 -278 1483 -273
rect 1510 -277 1512 -273
rect 1605 -278 1607 -273
rect 1620 -278 1622 -273
rect 1649 -277 1651 -273
rect 1729 -278 1731 -273
rect 1744 -278 1746 -273
rect 1773 -277 1775 -273
rect 682 -417 684 -412
rect 697 -417 699 -412
rect 726 -416 728 -412
rect 820 -417 822 -412
rect 835 -417 837 -412
rect 864 -416 866 -412
rect 966 -417 968 -412
rect 981 -417 983 -412
rect 1010 -416 1012 -412
rect 1090 -417 1092 -412
rect 1105 -417 1107 -412
rect 1134 -416 1136 -412
rect 1315 -417 1317 -412
rect 1330 -417 1332 -412
rect 1359 -416 1361 -412
rect 1462 -417 1464 -412
rect 1477 -417 1479 -412
rect 1506 -416 1508 -412
rect 1601 -417 1603 -412
rect 1616 -417 1618 -412
rect 1645 -416 1647 -412
rect 1725 -417 1727 -412
rect 1740 -417 1742 -412
rect 1769 -416 1771 -412
rect 1841 -461 1843 -456
rect 1856 -461 1858 -456
rect 1885 -460 1887 -456
rect 1841 -566 1843 -561
rect 1856 -566 1858 -561
rect 1885 -565 1887 -561
rect 3350 430 3352 440
rect 3365 430 3367 440
rect 3385 430 3387 440
rect 3395 430 3397 440
rect 3421 430 3423 440
rect 3668 480 3670 487
rect 3680 480 3682 487
rect 3695 480 3697 487
rect 3705 480 3707 487
rect 3728 480 3730 487
rect 2975 410 2977 414
rect 2978 343 2980 347
rect 2978 276 2980 280
rect 2996 171 2998 175
rect 2896 134 2898 139
rect 2915 134 2917 139
rect 2940 134 2942 139
rect 2959 134 2961 139
rect 2998 10 3000 14
rect 2898 -27 2900 -22
rect 2917 -27 2919 -22
rect 2942 -27 2944 -22
rect 2961 -27 2963 -22
rect 3488 392 3490 402
rect 3503 392 3505 402
rect 3523 392 3525 402
rect 3547 392 3549 402
rect 3614 352 3616 357
rect 3635 352 3637 357
rect 3661 353 3663 357
rect 3597 -44 3599 -34
rect 3612 -44 3614 -34
rect 3632 -44 3634 -34
rect 3642 -44 3644 -34
rect 3668 -44 3670 -34
rect 3709 -46 3711 -41
rect 3735 -46 3737 -41
rect 3767 -45 3769 -41
rect 2997 -144 2999 -140
rect 2897 -181 2899 -176
rect 2916 -181 2918 -176
rect 2941 -181 2943 -176
rect 2960 -181 2962 -176
rect 2997 -292 2999 -288
rect 3659 -300 3661 -293
rect 3671 -300 3673 -293
rect 3686 -300 3688 -293
rect 3696 -300 3698 -293
rect 3719 -300 3721 -293
rect 2897 -329 2899 -324
rect 2916 -329 2918 -324
rect 2941 -329 2943 -324
rect 2960 -329 2962 -324
rect 3434 -359 3436 -349
rect 3449 -359 3451 -349
rect 3464 -359 3466 -349
rect 3479 -359 3481 -349
rect 3493 -359 3495 -349
rect 3519 -359 3521 -349
rect 2973 -419 2975 -415
rect 3302 -443 3304 -433
rect 3317 -443 3319 -433
rect 3337 -443 3339 -433
rect 3347 -443 3349 -433
rect 3373 -443 3375 -433
rect 2975 -485 2977 -481
rect 3161 -518 3163 -508
rect 3176 -518 3178 -508
rect 3196 -518 3198 -508
rect 3220 -518 3222 -508
rect 2978 -552 2980 -548
rect 3063 -592 3065 -587
rect 3084 -592 3086 -587
rect 3110 -591 3112 -587
rect 2978 -619 2980 -615
rect 1841 -688 1843 -683
rect 1856 -688 1858 -683
rect 1885 -687 1887 -683
rect 1841 -795 1843 -790
rect 1856 -795 1858 -790
rect 1885 -794 1887 -790
<< ndiffusion >>
rect 2093 904 2098 905
rect 2097 900 2098 904
rect 2100 904 2104 905
rect 2112 904 2117 905
rect 2100 900 2102 904
rect 2116 900 2117 904
rect 2119 904 2125 905
rect 2119 900 2121 904
rect 2137 904 2142 905
rect 2141 900 2142 904
rect 2144 904 2150 905
rect 2144 900 2146 904
rect 2156 904 2161 905
rect 2160 900 2161 904
rect 2163 904 2169 905
rect 2163 900 2165 904
rect 2230 900 2235 901
rect 2234 896 2235 900
rect 2237 900 2241 901
rect 2249 900 2254 901
rect 2237 896 2239 900
rect 2253 896 2254 900
rect 2256 900 2262 901
rect 2256 896 2258 900
rect 2274 900 2279 901
rect 2278 896 2279 900
rect 2281 900 2287 901
rect 2281 896 2283 900
rect 2293 900 2298 901
rect 2297 896 2298 900
rect 2300 900 2306 901
rect 2300 896 2302 900
rect 2172 836 2173 840
rect 2175 836 2176 840
rect 2127 832 2129 836
rect 2123 829 2129 832
rect 2131 829 2144 836
rect 2146 833 2153 836
rect 2146 829 2149 833
rect 2392 845 2393 849
rect 2395 845 2396 849
rect 2345 835 2353 840
rect 2349 831 2353 835
rect 2355 836 2357 840
rect 2361 836 2362 840
rect 2355 831 2362 836
rect 2364 835 2372 840
rect 2364 831 2368 835
rect 2274 826 2275 830
rect 2277 826 2278 830
rect 2229 822 2231 826
rect 2225 819 2231 822
rect 2233 819 2246 826
rect 2248 823 2255 826
rect 2248 819 2251 823
rect 2091 628 2096 629
rect 2095 624 2096 628
rect 2098 628 2102 629
rect 2110 628 2115 629
rect 2098 624 2100 628
rect 2114 624 2115 628
rect 2117 628 2123 629
rect 2117 624 2119 628
rect 2135 628 2140 629
rect 2139 624 2140 628
rect 2142 628 2148 629
rect 2142 624 2144 628
rect 2154 628 2159 629
rect 2158 624 2159 628
rect 2161 628 2167 629
rect 2161 624 2163 628
rect 2228 624 2233 625
rect 2232 620 2233 624
rect 2235 624 2239 625
rect 2247 624 2252 625
rect 2235 620 2237 624
rect 2251 620 2252 624
rect 2254 624 2260 625
rect 2254 620 2256 624
rect 2272 624 2277 625
rect 2276 620 2277 624
rect 2279 624 2285 625
rect 2279 620 2281 624
rect 2291 624 2296 625
rect 2295 620 2296 624
rect 2298 624 2304 625
rect 2298 620 2300 624
rect 2170 560 2171 564
rect 2173 560 2174 564
rect 2125 556 2127 560
rect 2121 553 2127 556
rect 2129 553 2142 560
rect 2144 557 2151 560
rect 2144 553 2147 557
rect 2390 569 2391 573
rect 2393 569 2394 573
rect 2343 559 2351 564
rect 2347 555 2351 559
rect 2353 560 2355 564
rect 2359 560 2360 564
rect 2353 555 2360 560
rect 2362 559 2370 564
rect 2362 555 2366 559
rect 2272 550 2273 554
rect 2275 550 2276 554
rect 2227 546 2229 550
rect 2223 543 2229 546
rect 2231 543 2244 550
rect 2246 547 2253 550
rect 2246 543 2249 547
rect 2088 349 2093 350
rect 2092 345 2093 349
rect 2095 349 2099 350
rect 2107 349 2112 350
rect 2095 345 2097 349
rect 2111 345 2112 349
rect 2114 349 2120 350
rect 2114 345 2116 349
rect 2132 349 2137 350
rect 2136 345 2137 349
rect 2139 349 2145 350
rect 2139 345 2141 349
rect 2151 349 2156 350
rect 2155 345 2156 349
rect 2158 349 2164 350
rect 2158 345 2160 349
rect 2225 345 2230 346
rect 2229 341 2230 345
rect 2232 345 2236 346
rect 2244 345 2249 346
rect 2232 341 2234 345
rect 2248 341 2249 345
rect 2251 345 2257 346
rect 2251 341 2253 345
rect 2269 345 2274 346
rect 2273 341 2274 345
rect 2276 345 2282 346
rect 2276 341 2278 345
rect 2288 345 2293 346
rect 2292 341 2293 345
rect 2295 345 2301 346
rect 2295 341 2297 345
rect 2167 281 2168 285
rect 2170 281 2171 285
rect 2122 277 2124 281
rect 2118 274 2124 277
rect 2126 274 2139 281
rect 2141 278 2148 281
rect 2141 274 2144 278
rect 2387 290 2388 294
rect 2390 290 2391 294
rect 2340 280 2348 285
rect 2344 276 2348 280
rect 2350 281 2352 285
rect 2356 281 2357 285
rect 2350 276 2357 281
rect 2359 280 2367 285
rect 2359 276 2363 280
rect 2269 271 2270 275
rect 2272 271 2273 275
rect 2224 267 2226 271
rect 2220 264 2226 267
rect 2228 264 2241 271
rect 2243 268 2250 271
rect 2243 264 2246 268
rect 1428 3 1433 4
rect 1432 -1 1433 3
rect 1435 3 1439 4
rect 1447 3 1452 4
rect 1435 -1 1437 3
rect 1451 -1 1452 3
rect 1454 3 1460 4
rect 1454 -1 1456 3
rect 1472 3 1477 4
rect 1476 -1 1477 3
rect 1479 3 1485 4
rect 1479 -1 1481 3
rect 1491 3 1496 4
rect 1495 -1 1496 3
rect 1498 3 1504 4
rect 1498 -1 1500 3
rect 1577 1 1582 2
rect 1581 -3 1582 1
rect 1584 1 1588 2
rect 1596 1 1601 2
rect 1584 -3 1586 1
rect 1600 -3 1601 1
rect 1603 1 1609 2
rect 1603 -3 1605 1
rect 1621 1 1626 2
rect 1625 -3 1626 1
rect 1628 1 1634 2
rect 1628 -3 1630 1
rect 1640 1 1645 2
rect 1644 -3 1645 1
rect 1647 1 1653 2
rect 1647 -3 1649 1
rect 1729 0 1734 1
rect 1733 -4 1734 0
rect 1736 0 1740 1
rect 1748 0 1753 1
rect 1736 -4 1738 0
rect 1752 -4 1753 0
rect 1755 0 1761 1
rect 1755 -4 1757 0
rect 1773 0 1778 1
rect 1777 -4 1778 0
rect 1780 0 1786 1
rect 1780 -4 1782 0
rect 1792 0 1797 1
rect 1796 -4 1797 0
rect 1799 0 1805 1
rect 1799 -4 1801 0
rect 2091 64 2096 65
rect 2095 60 2096 64
rect 2098 64 2102 65
rect 2110 64 2115 65
rect 2098 60 2100 64
rect 2114 60 2115 64
rect 2117 64 2123 65
rect 2117 60 2119 64
rect 2135 64 2140 65
rect 2139 60 2140 64
rect 2142 64 2148 65
rect 2142 60 2144 64
rect 2154 64 2159 65
rect 2158 60 2159 64
rect 2161 64 2167 65
rect 2161 60 2163 64
rect 2228 60 2233 61
rect 2232 56 2233 60
rect 2235 60 2239 61
rect 2247 60 2252 61
rect 2235 56 2237 60
rect 2251 56 2252 60
rect 2254 60 2260 61
rect 2254 56 2256 60
rect 2272 60 2277 61
rect 2276 56 2277 60
rect 2279 60 2285 61
rect 2279 56 2281 60
rect 2291 60 2296 61
rect 2295 56 2296 60
rect 2298 60 2304 61
rect 2298 56 2300 60
rect 1880 -1 1885 0
rect 1884 -5 1885 -1
rect 1887 -1 1891 0
rect 1899 -1 1904 0
rect 1887 -5 1889 -1
rect 1903 -5 1904 -1
rect 1906 -1 1912 0
rect 1906 -5 1908 -1
rect 1924 -1 1929 0
rect 1928 -5 1929 -1
rect 1931 -1 1937 0
rect 1931 -5 1933 -1
rect 1943 -1 1948 0
rect 1947 -5 1948 -1
rect 1950 -1 1956 0
rect 1950 -5 1952 -1
rect 2170 -4 2171 0
rect 2173 -4 2174 0
rect 2125 -8 2127 -4
rect 2121 -11 2127 -8
rect 2129 -11 2142 -4
rect 2144 -7 2151 -4
rect 2144 -11 2147 -7
rect 2390 5 2391 9
rect 2393 5 2394 9
rect 2343 -5 2351 0
rect 2347 -9 2351 -5
rect 2353 -4 2355 0
rect 2359 -4 2360 0
rect 2353 -9 2360 -4
rect 2362 -5 2370 0
rect 2362 -9 2366 -5
rect 2272 -14 2273 -10
rect 2275 -14 2276 -10
rect 2227 -18 2229 -14
rect 2223 -21 2229 -18
rect 2231 -21 2244 -14
rect 2246 -17 2253 -14
rect 2246 -21 2249 -17
rect 109 -123 110 -119
rect 112 -123 113 -119
rect 430 -146 431 -142
rect 433 -146 434 -142
rect 376 -150 378 -146
rect 372 -153 378 -150
rect 380 -150 383 -146
rect 380 -153 387 -150
rect 402 -150 404 -146
rect 398 -153 404 -150
rect 406 -149 413 -146
rect 406 -153 409 -149
rect 1249 -84 1250 -80
rect 1252 -84 1253 -80
rect 1204 -88 1206 -84
rect 1200 -91 1206 -88
rect 1208 -91 1221 -84
rect 1223 -87 1230 -84
rect 1223 -91 1226 -87
rect 584 -168 585 -164
rect 587 -168 588 -164
rect 734 -168 735 -164
rect 737 -168 738 -164
rect 872 -168 873 -164
rect 875 -168 876 -164
rect 1018 -168 1019 -164
rect 1021 -168 1022 -164
rect 1142 -168 1143 -164
rect 1145 -168 1146 -164
rect 1367 -168 1368 -164
rect 1370 -168 1371 -164
rect 1514 -168 1515 -164
rect 1517 -168 1518 -164
rect 1653 -168 1654 -164
rect 1656 -168 1657 -164
rect 1777 -168 1778 -164
rect 1780 -168 1781 -164
rect 689 -172 691 -168
rect 109 -178 110 -174
rect 112 -178 113 -174
rect 537 -178 545 -173
rect 541 -182 545 -178
rect 547 -177 549 -173
rect 553 -177 554 -173
rect 547 -182 554 -177
rect 556 -178 564 -173
rect 685 -175 691 -172
rect 693 -175 706 -168
rect 708 -171 715 -168
rect 708 -175 711 -171
rect 827 -172 829 -168
rect 823 -175 829 -172
rect 831 -175 844 -168
rect 846 -171 853 -168
rect 846 -175 849 -171
rect 973 -172 975 -168
rect 969 -175 975 -172
rect 977 -175 990 -168
rect 992 -171 999 -168
rect 992 -175 995 -171
rect 1097 -172 1099 -168
rect 1093 -175 1099 -172
rect 1101 -175 1114 -168
rect 1116 -171 1123 -168
rect 1116 -175 1119 -171
rect 1322 -172 1324 -168
rect 1318 -175 1324 -172
rect 1326 -175 1339 -168
rect 1341 -171 1348 -168
rect 1341 -175 1344 -171
rect 1469 -172 1471 -168
rect 1465 -175 1471 -172
rect 1473 -175 1486 -168
rect 1488 -171 1495 -168
rect 1488 -175 1491 -171
rect 1608 -172 1610 -168
rect 1604 -175 1610 -172
rect 1612 -175 1625 -168
rect 1627 -171 1634 -168
rect 1627 -175 1630 -171
rect 1732 -172 1734 -168
rect 1728 -175 1734 -172
rect 1736 -175 1749 -168
rect 1751 -171 1758 -168
rect 1751 -175 1754 -171
rect 556 -182 560 -178
rect 430 -215 431 -211
rect 433 -215 434 -211
rect 376 -219 378 -215
rect 372 -222 378 -219
rect 380 -219 383 -215
rect 380 -222 387 -219
rect 402 -219 404 -215
rect 398 -222 404 -219
rect 406 -218 413 -215
rect 406 -222 409 -218
rect 3210 499 3219 505
rect 3214 495 3219 499
rect 3221 495 3234 505
rect 3236 495 3249 505
rect 3251 495 3264 505
rect 3266 495 3278 505
rect 3280 499 3289 505
rect 3280 495 3285 499
rect 3295 499 3304 505
rect 3299 495 3304 499
rect 3306 501 3311 505
rect 3306 495 3315 501
rect 430 -281 431 -277
rect 433 -281 434 -277
rect 376 -285 378 -281
rect 372 -288 378 -285
rect 380 -285 383 -281
rect 380 -288 387 -285
rect 402 -285 404 -281
rect 398 -288 404 -285
rect 406 -284 413 -281
rect 406 -288 409 -284
rect 729 -301 730 -297
rect 732 -301 733 -297
rect 684 -305 686 -301
rect 680 -308 686 -305
rect 688 -308 701 -301
rect 703 -304 710 -301
rect 703 -308 706 -304
rect 430 -347 431 -343
rect 433 -347 434 -343
rect 376 -351 378 -347
rect 372 -354 378 -351
rect 380 -351 383 -347
rect 380 -354 387 -351
rect 402 -351 404 -347
rect 398 -354 404 -351
rect 406 -350 413 -347
rect 406 -354 409 -350
rect 867 -301 868 -297
rect 870 -301 871 -297
rect 822 -305 824 -301
rect 818 -308 824 -305
rect 826 -308 839 -301
rect 841 -304 848 -301
rect 841 -308 844 -304
rect 1013 -301 1014 -297
rect 1016 -301 1017 -297
rect 968 -305 970 -301
rect 964 -308 970 -305
rect 972 -308 985 -301
rect 987 -304 994 -301
rect 987 -308 990 -304
rect 1137 -301 1138 -297
rect 1140 -301 1141 -297
rect 1092 -305 1094 -301
rect 1088 -308 1094 -305
rect 1096 -308 1109 -301
rect 1111 -304 1118 -301
rect 1111 -308 1114 -304
rect 1362 -301 1363 -297
rect 1365 -301 1366 -297
rect 1317 -305 1319 -301
rect 1313 -308 1319 -305
rect 1321 -308 1334 -301
rect 1336 -304 1343 -301
rect 1336 -308 1339 -304
rect 1509 -301 1510 -297
rect 1512 -301 1513 -297
rect 1464 -305 1466 -301
rect 1460 -308 1466 -305
rect 1468 -308 1481 -301
rect 1483 -304 1490 -301
rect 1483 -308 1486 -304
rect 1648 -301 1649 -297
rect 1651 -301 1652 -297
rect 1603 -305 1605 -301
rect 1599 -308 1605 -305
rect 1607 -308 1620 -301
rect 1622 -304 1629 -301
rect 1622 -308 1625 -304
rect 1772 -301 1773 -297
rect 1775 -301 1776 -297
rect 1727 -305 1729 -301
rect 1723 -308 1729 -305
rect 1731 -308 1744 -301
rect 1746 -304 1753 -301
rect 1746 -308 1749 -304
rect 725 -440 726 -436
rect 728 -440 729 -436
rect 680 -444 682 -440
rect 676 -447 682 -444
rect 684 -447 697 -440
rect 699 -443 706 -440
rect 699 -447 702 -443
rect 863 -440 864 -436
rect 866 -440 867 -436
rect 1009 -440 1010 -436
rect 1012 -440 1013 -436
rect 1133 -440 1134 -436
rect 1136 -440 1137 -436
rect 1358 -440 1359 -436
rect 1361 -440 1362 -436
rect 818 -444 820 -440
rect 814 -447 820 -444
rect 822 -447 835 -440
rect 837 -443 844 -440
rect 837 -447 840 -443
rect 964 -444 966 -440
rect 960 -447 966 -444
rect 968 -447 981 -440
rect 983 -443 990 -440
rect 983 -447 986 -443
rect 1088 -444 1090 -440
rect 1084 -447 1090 -444
rect 1092 -447 1105 -440
rect 1107 -443 1114 -440
rect 1107 -447 1110 -443
rect 1313 -444 1315 -440
rect 1309 -447 1315 -444
rect 1317 -447 1330 -440
rect 1332 -443 1339 -440
rect 1332 -447 1335 -443
rect 1505 -440 1506 -436
rect 1508 -440 1509 -436
rect 1460 -444 1462 -440
rect 1456 -447 1462 -444
rect 1464 -447 1477 -440
rect 1479 -443 1486 -440
rect 1479 -447 1482 -443
rect 1644 -440 1645 -436
rect 1647 -440 1648 -436
rect 1599 -444 1601 -440
rect 1595 -447 1601 -444
rect 1603 -447 1616 -440
rect 1618 -443 1625 -440
rect 1618 -447 1621 -443
rect 1768 -440 1769 -436
rect 1771 -440 1772 -436
rect 1723 -444 1725 -440
rect 1719 -447 1725 -444
rect 1727 -447 1740 -440
rect 1742 -443 1749 -440
rect 1742 -447 1745 -443
rect 1884 -484 1885 -480
rect 1887 -484 1888 -480
rect 1839 -488 1841 -484
rect 1835 -491 1841 -488
rect 1843 -491 1856 -484
rect 1858 -487 1865 -484
rect 1858 -491 1861 -487
rect 2972 452 2973 456
rect 2975 452 2976 456
rect 3660 454 3668 457
rect 3664 450 3668 454
rect 3670 453 3673 457
rect 3677 453 3680 457
rect 3670 450 3680 453
rect 3682 454 3695 457
rect 3682 450 3686 454
rect 3690 450 3695 454
rect 3697 453 3699 457
rect 3703 453 3705 457
rect 3697 450 3705 453
rect 3707 453 3712 457
rect 3707 450 3716 453
rect 3724 453 3728 457
rect 3720 450 3728 453
rect 3730 453 3733 457
rect 3730 450 3737 453
rect 3341 399 3350 405
rect 3345 395 3350 399
rect 3352 395 3365 405
rect 3367 395 3385 405
rect 3387 395 3395 405
rect 3397 399 3407 405
rect 3397 395 3403 399
rect 3412 399 3421 405
rect 3416 395 3421 399
rect 3423 401 3428 405
rect 3423 395 3432 401
rect 2974 386 2975 390
rect 2977 386 2978 390
rect 2977 319 2978 323
rect 2980 319 2981 323
rect 2977 252 2978 256
rect 2980 252 2981 256
rect 2995 147 2996 151
rect 2998 147 2999 151
rect 2891 107 2896 108
rect 2895 103 2896 107
rect 2898 107 2902 108
rect 2910 107 2915 108
rect 2898 103 2900 107
rect 2914 103 2915 107
rect 2917 107 2923 108
rect 2917 103 2919 107
rect 2935 107 2940 108
rect 2939 103 2940 107
rect 2942 107 2948 108
rect 2942 103 2944 107
rect 2954 107 2959 108
rect 2958 103 2959 107
rect 2961 107 2967 108
rect 2961 103 2963 107
rect 2997 -14 2998 -10
rect 3000 -14 3001 -10
rect 2893 -54 2898 -53
rect 2897 -58 2898 -54
rect 2900 -54 2904 -53
rect 2912 -54 2917 -53
rect 2900 -58 2902 -54
rect 2916 -58 2917 -54
rect 2919 -54 2925 -53
rect 2919 -58 2921 -54
rect 2937 -54 2942 -53
rect 2941 -58 2942 -54
rect 2944 -54 2950 -53
rect 2944 -58 2946 -54
rect 2956 -54 2961 -53
rect 2960 -58 2961 -54
rect 2963 -54 2969 -53
rect 2963 -58 2965 -54
rect 3479 361 3488 367
rect 3483 357 3488 361
rect 3490 357 3503 367
rect 3505 357 3523 367
rect 3525 361 3533 367
rect 3525 357 3529 361
rect 3538 361 3547 367
rect 3542 357 3547 361
rect 3549 363 3554 367
rect 3549 357 3558 363
rect 3660 329 3661 333
rect 3663 329 3664 333
rect 3612 325 3614 329
rect 3608 322 3614 325
rect 3616 322 3635 329
rect 3637 326 3644 329
rect 3637 322 3640 326
rect 3766 -69 3767 -65
rect 3769 -69 3770 -65
rect 3588 -75 3597 -69
rect 3592 -79 3597 -75
rect 3599 -79 3612 -69
rect 3614 -79 3632 -69
rect 3634 -79 3642 -69
rect 3644 -75 3654 -69
rect 3644 -79 3650 -75
rect 3659 -75 3668 -69
rect 3663 -79 3668 -75
rect 3670 -73 3675 -69
rect 3670 -79 3679 -73
rect 3707 -73 3709 -69
rect 3703 -76 3709 -73
rect 3711 -76 3735 -69
rect 3737 -72 3744 -69
rect 3737 -76 3740 -72
rect 2996 -168 2997 -164
rect 2999 -168 3000 -164
rect 2892 -208 2897 -207
rect 2896 -212 2897 -208
rect 2899 -208 2903 -207
rect 2911 -208 2916 -207
rect 2899 -212 2901 -208
rect 2915 -212 2916 -208
rect 2918 -208 2924 -207
rect 2918 -212 2920 -208
rect 2936 -208 2941 -207
rect 2940 -212 2941 -208
rect 2943 -208 2949 -207
rect 2943 -212 2945 -208
rect 2955 -208 2960 -207
rect 2959 -212 2960 -208
rect 2962 -208 2968 -207
rect 2962 -212 2964 -208
rect 2996 -316 2997 -312
rect 2999 -316 3000 -312
rect 3651 -326 3659 -323
rect 3655 -330 3659 -326
rect 3661 -327 3664 -323
rect 3668 -327 3671 -323
rect 3661 -330 3671 -327
rect 3673 -326 3686 -323
rect 3673 -330 3677 -326
rect 3681 -330 3686 -326
rect 3688 -327 3690 -323
rect 3694 -327 3696 -323
rect 3688 -330 3696 -327
rect 3698 -327 3703 -323
rect 3698 -330 3707 -327
rect 3715 -327 3719 -323
rect 3711 -330 3719 -327
rect 3721 -327 3724 -323
rect 3721 -330 3728 -327
rect 2892 -356 2897 -355
rect 2896 -360 2897 -356
rect 2899 -356 2903 -355
rect 2911 -356 2916 -355
rect 2899 -360 2901 -356
rect 2915 -360 2916 -356
rect 2918 -356 2924 -355
rect 2918 -360 2920 -356
rect 2936 -356 2941 -355
rect 2940 -360 2941 -356
rect 2943 -356 2949 -355
rect 2943 -360 2945 -356
rect 2955 -356 2960 -355
rect 2959 -360 2960 -356
rect 2962 -356 2968 -355
rect 2962 -360 2964 -356
rect 3425 -390 3434 -384
rect 3429 -394 3434 -390
rect 3436 -394 3449 -384
rect 3451 -394 3464 -384
rect 3466 -394 3479 -384
rect 3481 -394 3493 -384
rect 3495 -390 3504 -384
rect 3495 -394 3500 -390
rect 3510 -390 3519 -384
rect 3514 -394 3519 -390
rect 3521 -388 3526 -384
rect 3521 -394 3530 -388
rect 2972 -443 2973 -439
rect 2975 -443 2976 -439
rect 3293 -474 3302 -468
rect 3297 -478 3302 -474
rect 3304 -478 3317 -468
rect 3319 -478 3337 -468
rect 3339 -478 3347 -468
rect 3349 -474 3359 -468
rect 3349 -478 3355 -474
rect 3364 -474 3373 -468
rect 3368 -478 3373 -474
rect 3375 -472 3380 -468
rect 3375 -478 3384 -472
rect 2974 -509 2975 -505
rect 2977 -509 2978 -505
rect 3152 -549 3161 -543
rect 3156 -553 3161 -549
rect 3163 -553 3176 -543
rect 3178 -553 3196 -543
rect 3198 -549 3206 -543
rect 3198 -553 3202 -549
rect 3211 -549 3220 -543
rect 3215 -553 3220 -549
rect 3222 -547 3227 -543
rect 3222 -553 3231 -547
rect 2977 -576 2978 -572
rect 2980 -576 2981 -572
rect 1884 -589 1885 -585
rect 1887 -589 1888 -585
rect 1839 -593 1841 -589
rect 1835 -596 1841 -593
rect 1843 -596 1856 -589
rect 1858 -592 1865 -589
rect 1858 -596 1861 -592
rect 3109 -615 3110 -611
rect 3112 -615 3113 -611
rect 3061 -619 3063 -615
rect 3057 -622 3063 -619
rect 3065 -622 3084 -615
rect 3086 -618 3093 -615
rect 3086 -622 3089 -618
rect 2977 -643 2978 -639
rect 2980 -643 2981 -639
rect 1884 -711 1885 -707
rect 1887 -711 1888 -707
rect 1839 -715 1841 -711
rect 1835 -718 1841 -715
rect 1843 -718 1856 -711
rect 1858 -714 1865 -711
rect 1858 -718 1861 -714
rect 1884 -818 1885 -814
rect 1887 -818 1888 -814
rect 1839 -822 1841 -818
rect 1835 -825 1841 -822
rect 1843 -825 1856 -818
rect 1858 -821 1865 -818
rect 1858 -825 1861 -821
<< pdiffusion >>
rect 2093 935 2098 936
rect 2097 931 2098 935
rect 2100 935 2106 936
rect 2100 931 2102 935
rect 2112 935 2117 936
rect 2116 931 2117 935
rect 2119 935 2125 936
rect 2119 931 2121 935
rect 2137 935 2142 936
rect 2141 931 2142 935
rect 2144 935 2150 936
rect 2144 931 2146 935
rect 2156 935 2161 936
rect 2160 931 2161 935
rect 2163 935 2169 936
rect 2163 931 2165 935
rect 2230 931 2235 932
rect 2234 927 2235 931
rect 2237 931 2243 932
rect 2237 927 2239 931
rect 2249 931 2254 932
rect 2253 927 2254 931
rect 2256 931 2262 932
rect 2256 927 2258 931
rect 2274 931 2279 932
rect 2278 927 2279 931
rect 2281 931 2287 932
rect 2281 927 2283 931
rect 2293 931 2298 932
rect 2297 927 2298 931
rect 2300 931 2306 932
rect 2300 927 2302 931
rect 2349 869 2353 873
rect 2345 864 2353 869
rect 2355 864 2362 873
rect 2364 868 2372 873
rect 2392 869 2393 873
rect 2395 869 2396 873
rect 2364 864 2368 868
rect 2123 863 2129 864
rect 2127 859 2129 863
rect 2131 860 2135 864
rect 2139 860 2144 864
rect 2131 859 2144 860
rect 2146 863 2153 864
rect 2146 859 2149 863
rect 2172 860 2173 864
rect 2175 860 2176 864
rect 2225 853 2231 854
rect 2229 849 2231 853
rect 2233 850 2237 854
rect 2241 850 2246 854
rect 2233 849 2246 850
rect 2248 853 2255 854
rect 2248 849 2251 853
rect 2274 850 2275 854
rect 2277 850 2278 854
rect 2091 659 2096 660
rect 2095 655 2096 659
rect 2098 659 2104 660
rect 2098 655 2100 659
rect 2110 659 2115 660
rect 2114 655 2115 659
rect 2117 659 2123 660
rect 2117 655 2119 659
rect 2135 659 2140 660
rect 2139 655 2140 659
rect 2142 659 2148 660
rect 2142 655 2144 659
rect 2154 659 2159 660
rect 2158 655 2159 659
rect 2161 659 2167 660
rect 2161 655 2163 659
rect 2228 655 2233 656
rect 2232 651 2233 655
rect 2235 655 2241 656
rect 2235 651 2237 655
rect 2247 655 2252 656
rect 2251 651 2252 655
rect 2254 655 2260 656
rect 2254 651 2256 655
rect 2272 655 2277 656
rect 2276 651 2277 655
rect 2279 655 2285 656
rect 2279 651 2281 655
rect 2291 655 2296 656
rect 2295 651 2296 655
rect 2298 655 2304 656
rect 2298 651 2300 655
rect 2347 593 2351 597
rect 2343 588 2351 593
rect 2353 588 2360 597
rect 2362 592 2370 597
rect 2390 593 2391 597
rect 2393 593 2394 597
rect 2362 588 2366 592
rect 2121 587 2127 588
rect 2125 583 2127 587
rect 2129 584 2133 588
rect 2137 584 2142 588
rect 2129 583 2142 584
rect 2144 587 2151 588
rect 2144 583 2147 587
rect 2170 584 2171 588
rect 2173 584 2174 588
rect 2223 577 2229 578
rect 2227 573 2229 577
rect 2231 574 2235 578
rect 2239 574 2244 578
rect 2231 573 2244 574
rect 2246 577 2253 578
rect 2246 573 2249 577
rect 2272 574 2273 578
rect 2275 574 2276 578
rect 2088 380 2093 381
rect 2092 376 2093 380
rect 2095 380 2101 381
rect 2095 376 2097 380
rect 2107 380 2112 381
rect 2111 376 2112 380
rect 2114 380 2120 381
rect 2114 376 2116 380
rect 2132 380 2137 381
rect 2136 376 2137 380
rect 2139 380 2145 381
rect 2139 376 2141 380
rect 2151 380 2156 381
rect 2155 376 2156 380
rect 2158 380 2164 381
rect 2158 376 2160 380
rect 2225 376 2230 377
rect 2229 372 2230 376
rect 2232 376 2238 377
rect 2232 372 2234 376
rect 2244 376 2249 377
rect 2248 372 2249 376
rect 2251 376 2257 377
rect 2251 372 2253 376
rect 2269 376 2274 377
rect 2273 372 2274 376
rect 2276 376 2282 377
rect 2276 372 2278 376
rect 2288 376 2293 377
rect 2292 372 2293 376
rect 2295 376 2301 377
rect 2295 372 2297 376
rect 2344 314 2348 318
rect 2340 309 2348 314
rect 2350 309 2357 318
rect 2359 313 2367 318
rect 2387 314 2388 318
rect 2390 314 2391 318
rect 2359 309 2363 313
rect 2118 308 2124 309
rect 2122 304 2124 308
rect 2126 305 2130 309
rect 2134 305 2139 309
rect 2126 304 2139 305
rect 2141 308 2148 309
rect 2141 304 2144 308
rect 2167 305 2168 309
rect 2170 305 2171 309
rect 2220 298 2226 299
rect 2224 294 2226 298
rect 2228 295 2232 299
rect 2236 295 2241 299
rect 2228 294 2241 295
rect 2243 298 2250 299
rect 2243 294 2246 298
rect 2269 295 2270 299
rect 2272 295 2273 299
rect 1428 34 1433 35
rect 1432 30 1433 34
rect 1435 34 1441 35
rect 1435 30 1437 34
rect 1447 34 1452 35
rect 1451 30 1452 34
rect 1454 34 1460 35
rect 1454 30 1456 34
rect 1472 34 1477 35
rect 1476 30 1477 34
rect 1479 34 1485 35
rect 1479 30 1481 34
rect 1491 34 1496 35
rect 1495 30 1496 34
rect 1498 34 1504 35
rect 1498 30 1500 34
rect 1577 32 1582 33
rect 1581 28 1582 32
rect 1584 32 1590 33
rect 1584 28 1586 32
rect 1596 32 1601 33
rect 1600 28 1601 32
rect 1603 32 1609 33
rect 1603 28 1605 32
rect 1621 32 1626 33
rect 1625 28 1626 32
rect 1628 32 1634 33
rect 1628 28 1630 32
rect 1640 32 1645 33
rect 1644 28 1645 32
rect 1647 32 1653 33
rect 1647 28 1649 32
rect 1729 31 1734 32
rect 1733 27 1734 31
rect 1736 31 1742 32
rect 1736 27 1738 31
rect 1748 31 1753 32
rect 1752 27 1753 31
rect 1755 31 1761 32
rect 1755 27 1757 31
rect 1773 31 1778 32
rect 1777 27 1778 31
rect 1780 31 1786 32
rect 1780 27 1782 31
rect 1792 31 1797 32
rect 1796 27 1797 31
rect 1799 31 1805 32
rect 1799 27 1801 31
rect 2091 95 2096 96
rect 2095 91 2096 95
rect 2098 95 2104 96
rect 2098 91 2100 95
rect 2110 95 2115 96
rect 2114 91 2115 95
rect 2117 95 2123 96
rect 2117 91 2119 95
rect 2135 95 2140 96
rect 2139 91 2140 95
rect 2142 95 2148 96
rect 2142 91 2144 95
rect 2154 95 2159 96
rect 2158 91 2159 95
rect 2161 95 2167 96
rect 2161 91 2163 95
rect 2228 91 2233 92
rect 2232 87 2233 91
rect 2235 91 2241 92
rect 2235 87 2237 91
rect 2247 91 2252 92
rect 2251 87 2252 91
rect 2254 91 2260 92
rect 2254 87 2256 91
rect 2272 91 2277 92
rect 2276 87 2277 91
rect 2279 91 2285 92
rect 2279 87 2281 91
rect 2291 91 2296 92
rect 2295 87 2296 91
rect 2298 91 2304 92
rect 2298 87 2300 91
rect 1880 30 1885 31
rect 1884 26 1885 30
rect 1887 30 1893 31
rect 1887 26 1889 30
rect 1899 30 1904 31
rect 1903 26 1904 30
rect 1906 30 1912 31
rect 1906 26 1908 30
rect 1924 30 1929 31
rect 1928 26 1929 30
rect 1931 30 1937 31
rect 1931 26 1933 30
rect 1943 30 1948 31
rect 1947 26 1948 30
rect 1950 30 1956 31
rect 1950 26 1952 30
rect 2347 29 2351 33
rect 2343 24 2351 29
rect 2353 24 2360 33
rect 2362 28 2370 33
rect 2390 29 2391 33
rect 2393 29 2394 33
rect 2362 24 2366 28
rect 2121 23 2127 24
rect 2125 19 2127 23
rect 2129 20 2133 24
rect 2137 20 2142 24
rect 2129 19 2142 20
rect 2144 23 2151 24
rect 2144 19 2147 23
rect 2170 20 2171 24
rect 2173 20 2174 24
rect 2223 13 2229 14
rect 2227 9 2229 13
rect 2231 10 2235 14
rect 2239 10 2244 14
rect 2231 9 2244 10
rect 2246 13 2253 14
rect 2246 9 2249 13
rect 2272 10 2273 14
rect 2275 10 2276 14
rect 1200 -57 1206 -56
rect 1204 -61 1206 -57
rect 1208 -60 1212 -56
rect 1216 -60 1221 -56
rect 1208 -61 1221 -60
rect 1223 -57 1230 -56
rect 1223 -61 1226 -57
rect 1249 -60 1250 -56
rect 1252 -60 1253 -56
rect 109 -99 110 -95
rect 112 -99 113 -95
rect 372 -119 378 -118
rect 376 -123 378 -119
rect 380 -122 383 -118
rect 380 -123 387 -122
rect 398 -119 404 -118
rect 402 -123 404 -119
rect 406 -122 409 -118
rect 430 -122 431 -118
rect 433 -122 434 -118
rect 406 -123 413 -122
rect 109 -154 110 -150
rect 112 -154 113 -150
rect 541 -144 545 -140
rect 537 -149 545 -144
rect 547 -149 554 -140
rect 556 -145 564 -140
rect 584 -144 585 -140
rect 587 -144 588 -140
rect 556 -149 560 -145
rect 685 -141 691 -140
rect 689 -145 691 -141
rect 693 -144 697 -140
rect 701 -144 706 -140
rect 693 -145 706 -144
rect 708 -141 715 -140
rect 708 -145 711 -141
rect 734 -144 735 -140
rect 737 -144 738 -140
rect 823 -141 829 -140
rect 827 -145 829 -141
rect 831 -144 835 -140
rect 839 -144 844 -140
rect 831 -145 844 -144
rect 846 -141 853 -140
rect 846 -145 849 -141
rect 872 -144 873 -140
rect 875 -144 876 -140
rect 969 -141 975 -140
rect 973 -145 975 -141
rect 977 -144 981 -140
rect 985 -144 990 -140
rect 977 -145 990 -144
rect 992 -141 999 -140
rect 992 -145 995 -141
rect 1018 -144 1019 -140
rect 1021 -144 1022 -140
rect 1093 -141 1099 -140
rect 1097 -145 1099 -141
rect 1101 -144 1105 -140
rect 1109 -144 1114 -140
rect 1101 -145 1114 -144
rect 1116 -141 1123 -140
rect 1116 -145 1119 -141
rect 1142 -144 1143 -140
rect 1145 -144 1146 -140
rect 1318 -141 1324 -140
rect 1322 -145 1324 -141
rect 1326 -144 1330 -140
rect 1334 -144 1339 -140
rect 1326 -145 1339 -144
rect 1341 -141 1348 -140
rect 1341 -145 1344 -141
rect 1367 -144 1368 -140
rect 1370 -144 1371 -140
rect 1465 -141 1471 -140
rect 1469 -145 1471 -141
rect 1473 -144 1477 -140
rect 1481 -144 1486 -140
rect 1473 -145 1486 -144
rect 1488 -141 1495 -140
rect 1488 -145 1491 -141
rect 1514 -144 1515 -140
rect 1517 -144 1518 -140
rect 1604 -141 1610 -140
rect 1608 -145 1610 -141
rect 1612 -144 1616 -140
rect 1620 -144 1625 -140
rect 1612 -145 1625 -144
rect 1627 -141 1634 -140
rect 1627 -145 1630 -141
rect 1653 -144 1654 -140
rect 1656 -144 1657 -140
rect 1728 -141 1734 -140
rect 1732 -145 1734 -141
rect 1736 -144 1740 -140
rect 1744 -144 1749 -140
rect 1736 -145 1749 -144
rect 1751 -141 1758 -140
rect 1751 -145 1754 -141
rect 1777 -144 1778 -140
rect 1780 -144 1781 -140
rect 372 -188 378 -187
rect 376 -192 378 -188
rect 380 -191 383 -187
rect 380 -192 387 -191
rect 398 -188 404 -187
rect 402 -192 404 -188
rect 406 -191 409 -187
rect 430 -191 431 -187
rect 433 -191 434 -187
rect 406 -192 413 -191
rect 372 -254 378 -253
rect 376 -258 378 -254
rect 380 -257 383 -253
rect 380 -258 387 -257
rect 398 -254 404 -253
rect 402 -258 404 -254
rect 406 -257 409 -253
rect 430 -257 431 -253
rect 433 -257 434 -253
rect 3210 534 3219 540
rect 3214 530 3219 534
rect 3221 534 3234 540
rect 3221 530 3223 534
rect 3227 530 3234 534
rect 3236 534 3249 540
rect 3236 530 3240 534
rect 3244 530 3249 534
rect 3251 534 3264 540
rect 3251 530 3255 534
rect 3259 530 3264 534
rect 3266 534 3278 540
rect 3266 530 3270 534
rect 3274 530 3278 534
rect 3280 534 3289 540
rect 3280 530 3285 534
rect 3295 534 3304 540
rect 3299 530 3304 534
rect 3306 534 3315 540
rect 3306 530 3311 534
rect 2972 476 2973 480
rect 2975 476 2976 480
rect 406 -258 413 -257
rect 680 -274 686 -273
rect 684 -278 686 -274
rect 688 -277 692 -273
rect 696 -277 701 -273
rect 688 -278 701 -277
rect 703 -274 710 -273
rect 703 -278 706 -274
rect 729 -277 730 -273
rect 732 -277 733 -273
rect 818 -274 824 -273
rect 822 -278 824 -274
rect 826 -277 830 -273
rect 834 -277 839 -273
rect 826 -278 839 -277
rect 841 -274 848 -273
rect 841 -278 844 -274
rect 867 -277 868 -273
rect 870 -277 871 -273
rect 372 -320 378 -319
rect 376 -324 378 -320
rect 380 -323 383 -319
rect 380 -324 387 -323
rect 398 -320 404 -319
rect 402 -324 404 -320
rect 406 -323 409 -319
rect 430 -323 431 -319
rect 433 -323 434 -319
rect 406 -324 413 -323
rect 964 -274 970 -273
rect 968 -278 970 -274
rect 972 -277 976 -273
rect 980 -277 985 -273
rect 972 -278 985 -277
rect 987 -274 994 -273
rect 987 -278 990 -274
rect 1013 -277 1014 -273
rect 1016 -277 1017 -273
rect 1088 -274 1094 -273
rect 1092 -278 1094 -274
rect 1096 -277 1100 -273
rect 1104 -277 1109 -273
rect 1096 -278 1109 -277
rect 1111 -274 1118 -273
rect 1111 -278 1114 -274
rect 1137 -277 1138 -273
rect 1140 -277 1141 -273
rect 1313 -274 1319 -273
rect 1317 -278 1319 -274
rect 1321 -277 1325 -273
rect 1329 -277 1334 -273
rect 1321 -278 1334 -277
rect 1336 -274 1343 -273
rect 1336 -278 1339 -274
rect 1362 -277 1363 -273
rect 1365 -277 1366 -273
rect 1460 -274 1466 -273
rect 1464 -278 1466 -274
rect 1468 -277 1472 -273
rect 1476 -277 1481 -273
rect 1468 -278 1481 -277
rect 1483 -274 1490 -273
rect 1483 -278 1486 -274
rect 1509 -277 1510 -273
rect 1512 -277 1513 -273
rect 1599 -274 1605 -273
rect 1603 -278 1605 -274
rect 1607 -277 1611 -273
rect 1615 -277 1620 -273
rect 1607 -278 1620 -277
rect 1622 -274 1629 -273
rect 1622 -278 1625 -274
rect 1648 -277 1649 -273
rect 1651 -277 1652 -273
rect 1723 -274 1729 -273
rect 1727 -278 1729 -274
rect 1731 -277 1735 -273
rect 1739 -277 1744 -273
rect 1731 -278 1744 -277
rect 1746 -274 1753 -273
rect 1746 -278 1749 -274
rect 1772 -277 1773 -273
rect 1775 -277 1776 -273
rect 676 -413 682 -412
rect 680 -417 682 -413
rect 684 -416 688 -412
rect 692 -416 697 -412
rect 684 -417 697 -416
rect 699 -413 706 -412
rect 699 -417 702 -413
rect 725 -416 726 -412
rect 728 -416 729 -412
rect 814 -413 820 -412
rect 818 -417 820 -413
rect 822 -416 826 -412
rect 830 -416 835 -412
rect 822 -417 835 -416
rect 837 -413 844 -412
rect 837 -417 840 -413
rect 863 -416 864 -412
rect 866 -416 867 -412
rect 960 -413 966 -412
rect 964 -417 966 -413
rect 968 -416 972 -412
rect 976 -416 981 -412
rect 968 -417 981 -416
rect 983 -413 990 -412
rect 983 -417 986 -413
rect 1009 -416 1010 -412
rect 1012 -416 1013 -412
rect 1084 -413 1090 -412
rect 1088 -417 1090 -413
rect 1092 -416 1096 -412
rect 1100 -416 1105 -412
rect 1092 -417 1105 -416
rect 1107 -413 1114 -412
rect 1107 -417 1110 -413
rect 1133 -416 1134 -412
rect 1136 -416 1137 -412
rect 1309 -413 1315 -412
rect 1313 -417 1315 -413
rect 1317 -416 1321 -412
rect 1325 -416 1330 -412
rect 1317 -417 1330 -416
rect 1332 -413 1339 -412
rect 1332 -417 1335 -413
rect 1358 -416 1359 -412
rect 1361 -416 1362 -412
rect 1456 -413 1462 -412
rect 1460 -417 1462 -413
rect 1464 -416 1468 -412
rect 1472 -416 1477 -412
rect 1464 -417 1477 -416
rect 1479 -413 1486 -412
rect 1479 -417 1482 -413
rect 1505 -416 1506 -412
rect 1508 -416 1509 -412
rect 1595 -413 1601 -412
rect 1599 -417 1601 -413
rect 1603 -416 1607 -412
rect 1611 -416 1616 -412
rect 1603 -417 1616 -416
rect 1618 -413 1625 -412
rect 1618 -417 1621 -413
rect 1644 -416 1645 -412
rect 1647 -416 1648 -412
rect 1719 -413 1725 -412
rect 1723 -417 1725 -413
rect 1727 -416 1731 -412
rect 1735 -416 1740 -412
rect 1727 -417 1740 -416
rect 1742 -413 1749 -412
rect 1742 -417 1745 -413
rect 1768 -416 1769 -412
rect 1771 -416 1772 -412
rect 1835 -457 1841 -456
rect 1839 -461 1841 -457
rect 1843 -460 1847 -456
rect 1851 -460 1856 -456
rect 1843 -461 1856 -460
rect 1858 -457 1865 -456
rect 1858 -461 1861 -457
rect 1884 -460 1885 -456
rect 1887 -460 1888 -456
rect 1835 -562 1841 -561
rect 1839 -566 1841 -562
rect 1843 -565 1847 -561
rect 1851 -565 1856 -561
rect 1843 -566 1856 -565
rect 1858 -562 1865 -561
rect 1858 -566 1861 -562
rect 1884 -565 1885 -561
rect 1887 -565 1888 -561
rect 3341 434 3350 440
rect 3345 430 3350 434
rect 3352 434 3365 440
rect 3352 430 3356 434
rect 3361 430 3365 434
rect 3367 434 3385 440
rect 3367 430 3374 434
rect 3378 430 3385 434
rect 3387 434 3395 440
rect 3387 430 3389 434
rect 3393 430 3395 434
rect 3397 434 3407 440
rect 3397 430 3403 434
rect 3412 434 3421 440
rect 3416 430 3421 434
rect 3423 434 3432 440
rect 3423 430 3428 434
rect 3660 484 3668 487
rect 3664 480 3668 484
rect 3670 480 3680 487
rect 3682 480 3695 487
rect 3697 480 3705 487
rect 3707 484 3716 487
rect 3707 480 3712 484
rect 3720 484 3728 487
rect 3724 480 3728 484
rect 3730 484 3737 487
rect 3730 480 3733 484
rect 2974 410 2975 414
rect 2977 410 2978 414
rect 3479 396 3488 402
rect 2977 343 2978 347
rect 2980 343 2981 347
rect 2977 276 2978 280
rect 2980 276 2981 280
rect 2995 171 2996 175
rect 2998 171 2999 175
rect 2891 138 2896 139
rect 2895 134 2896 138
rect 2898 138 2904 139
rect 2898 134 2900 138
rect 2910 138 2915 139
rect 2914 134 2915 138
rect 2917 138 2923 139
rect 2917 134 2919 138
rect 2935 138 2940 139
rect 2939 134 2940 138
rect 2942 138 2948 139
rect 2942 134 2944 138
rect 2954 138 2959 139
rect 2958 134 2959 138
rect 2961 138 2967 139
rect 2961 134 2963 138
rect 2997 10 2998 14
rect 3000 10 3001 14
rect 2893 -23 2898 -22
rect 2897 -27 2898 -23
rect 2900 -23 2906 -22
rect 2900 -27 2902 -23
rect 2912 -23 2917 -22
rect 2916 -27 2917 -23
rect 2919 -23 2925 -22
rect 2919 -27 2921 -23
rect 2937 -23 2942 -22
rect 2941 -27 2942 -23
rect 2944 -23 2950 -22
rect 2944 -27 2946 -23
rect 2956 -23 2961 -22
rect 2960 -27 2961 -23
rect 2963 -23 2969 -22
rect 2963 -27 2965 -23
rect 3483 392 3488 396
rect 3490 396 3503 402
rect 3490 392 3494 396
rect 3499 392 3503 396
rect 3505 396 3523 402
rect 3505 392 3512 396
rect 3516 392 3523 396
rect 3525 396 3533 402
rect 3525 392 3529 396
rect 3538 396 3547 402
rect 3542 392 3547 396
rect 3549 396 3558 402
rect 3549 392 3554 396
rect 3608 356 3614 357
rect 3612 352 3614 356
rect 3616 353 3619 357
rect 3616 352 3623 353
rect 3629 356 3635 357
rect 3633 352 3635 356
rect 3637 353 3640 357
rect 3660 353 3661 357
rect 3663 353 3664 357
rect 3637 352 3644 353
rect 3588 -40 3597 -34
rect 3592 -44 3597 -40
rect 3599 -40 3612 -34
rect 3599 -44 3603 -40
rect 3608 -44 3612 -40
rect 3614 -40 3632 -34
rect 3614 -44 3621 -40
rect 3625 -44 3632 -40
rect 3634 -40 3642 -34
rect 3634 -44 3636 -40
rect 3640 -44 3642 -40
rect 3644 -40 3654 -34
rect 3644 -44 3650 -40
rect 3659 -40 3668 -34
rect 3663 -44 3668 -40
rect 3670 -40 3679 -34
rect 3670 -44 3675 -40
rect 3703 -42 3709 -41
rect 3707 -46 3709 -42
rect 3711 -45 3714 -41
rect 3711 -46 3718 -45
rect 3729 -42 3735 -41
rect 3733 -46 3735 -42
rect 3737 -45 3740 -41
rect 3766 -45 3767 -41
rect 3769 -45 3770 -41
rect 3737 -46 3744 -45
rect 2996 -144 2997 -140
rect 2999 -144 3000 -140
rect 2892 -177 2897 -176
rect 2896 -181 2897 -177
rect 2899 -177 2905 -176
rect 2899 -181 2901 -177
rect 2911 -177 2916 -176
rect 2915 -181 2916 -177
rect 2918 -177 2924 -176
rect 2918 -181 2920 -177
rect 2936 -177 2941 -176
rect 2940 -181 2941 -177
rect 2943 -177 2949 -176
rect 2943 -181 2945 -177
rect 2955 -177 2960 -176
rect 2959 -181 2960 -177
rect 2962 -177 2968 -176
rect 2962 -181 2964 -177
rect 2996 -292 2997 -288
rect 2999 -292 3000 -288
rect 3651 -296 3659 -293
rect 3655 -300 3659 -296
rect 3661 -300 3671 -293
rect 3673 -300 3686 -293
rect 3688 -300 3696 -293
rect 3698 -296 3707 -293
rect 3698 -300 3703 -296
rect 3711 -296 3719 -293
rect 3715 -300 3719 -296
rect 3721 -296 3728 -293
rect 3721 -300 3724 -296
rect 2892 -325 2897 -324
rect 2896 -329 2897 -325
rect 2899 -325 2905 -324
rect 2899 -329 2901 -325
rect 2911 -325 2916 -324
rect 2915 -329 2916 -325
rect 2918 -325 2924 -324
rect 2918 -329 2920 -325
rect 2936 -325 2941 -324
rect 2940 -329 2941 -325
rect 2943 -325 2949 -324
rect 2943 -329 2945 -325
rect 2955 -325 2960 -324
rect 2959 -329 2960 -325
rect 2962 -325 2968 -324
rect 2962 -329 2964 -325
rect 3425 -355 3434 -349
rect 3429 -359 3434 -355
rect 3436 -355 3449 -349
rect 3436 -359 3438 -355
rect 3442 -359 3449 -355
rect 3451 -355 3464 -349
rect 3451 -359 3455 -355
rect 3459 -359 3464 -355
rect 3466 -355 3479 -349
rect 3466 -359 3470 -355
rect 3474 -359 3479 -355
rect 3481 -355 3493 -349
rect 3481 -359 3485 -355
rect 3489 -359 3493 -355
rect 3495 -355 3504 -349
rect 3495 -359 3500 -355
rect 3510 -355 3519 -349
rect 3514 -359 3519 -355
rect 3521 -355 3530 -349
rect 3521 -359 3526 -355
rect 2972 -419 2973 -415
rect 2975 -419 2976 -415
rect 3293 -439 3302 -433
rect 3297 -443 3302 -439
rect 3304 -439 3317 -433
rect 3304 -443 3308 -439
rect 3313 -443 3317 -439
rect 3319 -439 3337 -433
rect 3319 -443 3326 -439
rect 3330 -443 3337 -439
rect 3339 -439 3347 -433
rect 3339 -443 3341 -439
rect 3345 -443 3347 -439
rect 3349 -439 3359 -433
rect 3349 -443 3355 -439
rect 3364 -439 3373 -433
rect 3368 -443 3373 -439
rect 3375 -439 3384 -433
rect 3375 -443 3380 -439
rect 2974 -485 2975 -481
rect 2977 -485 2978 -481
rect 3152 -514 3161 -508
rect 3156 -518 3161 -514
rect 3163 -514 3176 -508
rect 3163 -518 3167 -514
rect 3172 -518 3176 -514
rect 3178 -514 3196 -508
rect 3178 -518 3185 -514
rect 3189 -518 3196 -514
rect 3198 -514 3206 -508
rect 3198 -518 3202 -514
rect 3211 -514 3220 -508
rect 3215 -518 3220 -514
rect 3222 -514 3231 -508
rect 3222 -518 3227 -514
rect 2977 -552 2978 -548
rect 2980 -552 2981 -548
rect 3057 -588 3063 -587
rect 3061 -592 3063 -588
rect 3065 -591 3068 -587
rect 3065 -592 3072 -591
rect 3078 -588 3084 -587
rect 3082 -592 3084 -588
rect 3086 -591 3089 -587
rect 3109 -591 3110 -587
rect 3112 -591 3113 -587
rect 3086 -592 3093 -591
rect 2977 -619 2978 -615
rect 2980 -619 2981 -615
rect 1835 -684 1841 -683
rect 1839 -688 1841 -684
rect 1843 -687 1847 -683
rect 1851 -687 1856 -683
rect 1843 -688 1856 -687
rect 1858 -684 1865 -683
rect 1858 -688 1861 -684
rect 1884 -687 1885 -683
rect 1887 -687 1888 -683
rect 1835 -791 1841 -790
rect 1839 -795 1841 -791
rect 1843 -794 1847 -790
rect 1851 -794 1856 -790
rect 1843 -795 1856 -794
rect 1858 -791 1865 -790
rect 1858 -795 1861 -791
rect 1884 -794 1885 -790
rect 1887 -794 1888 -790
<< ndcontact >>
rect 2093 900 2097 904
rect 2102 900 2106 904
rect 2112 900 2116 904
rect 2121 900 2125 904
rect 2137 900 2141 904
rect 2146 900 2150 904
rect 2156 900 2160 904
rect 2165 900 2169 904
rect 2230 896 2234 900
rect 2239 896 2243 900
rect 2249 896 2253 900
rect 2258 896 2262 900
rect 2274 896 2278 900
rect 2283 896 2287 900
rect 2293 896 2297 900
rect 2302 896 2306 900
rect 2168 836 2172 840
rect 2176 836 2180 840
rect 2123 832 2127 836
rect 2149 829 2153 833
rect 2388 845 2392 849
rect 2396 845 2400 849
rect 2345 831 2349 835
rect 2357 836 2361 840
rect 2368 831 2372 835
rect 2270 826 2274 830
rect 2278 826 2282 830
rect 2225 822 2229 826
rect 2251 819 2255 823
rect 2091 624 2095 628
rect 2100 624 2104 628
rect 2110 624 2114 628
rect 2119 624 2123 628
rect 2135 624 2139 628
rect 2144 624 2148 628
rect 2154 624 2158 628
rect 2163 624 2167 628
rect 2228 620 2232 624
rect 2237 620 2241 624
rect 2247 620 2251 624
rect 2256 620 2260 624
rect 2272 620 2276 624
rect 2281 620 2285 624
rect 2291 620 2295 624
rect 2300 620 2304 624
rect 2166 560 2170 564
rect 2174 560 2178 564
rect 2121 556 2125 560
rect 2147 553 2151 557
rect 2386 569 2390 573
rect 2394 569 2398 573
rect 2343 555 2347 559
rect 2355 560 2359 564
rect 2366 555 2370 559
rect 2268 550 2272 554
rect 2276 550 2280 554
rect 2223 546 2227 550
rect 2249 543 2253 547
rect 2088 345 2092 349
rect 2097 345 2101 349
rect 2107 345 2111 349
rect 2116 345 2120 349
rect 2132 345 2136 349
rect 2141 345 2145 349
rect 2151 345 2155 349
rect 2160 345 2164 349
rect 2225 341 2229 345
rect 2234 341 2238 345
rect 2244 341 2248 345
rect 2253 341 2257 345
rect 2269 341 2273 345
rect 2278 341 2282 345
rect 2288 341 2292 345
rect 2297 341 2301 345
rect 2163 281 2167 285
rect 2171 281 2175 285
rect 2118 277 2122 281
rect 2144 274 2148 278
rect 2383 290 2387 294
rect 2391 290 2395 294
rect 2340 276 2344 280
rect 2352 281 2356 285
rect 2363 276 2367 280
rect 2265 271 2269 275
rect 2273 271 2277 275
rect 2220 267 2224 271
rect 2246 264 2250 268
rect 1428 -1 1432 3
rect 1437 -1 1441 3
rect 1447 -1 1451 3
rect 1456 -1 1460 3
rect 1472 -1 1476 3
rect 1481 -1 1485 3
rect 1491 -1 1495 3
rect 1500 -1 1504 3
rect 1577 -3 1581 1
rect 1586 -3 1590 1
rect 1596 -3 1600 1
rect 1605 -3 1609 1
rect 1621 -3 1625 1
rect 1630 -3 1634 1
rect 1640 -3 1644 1
rect 1649 -3 1653 1
rect 1729 -4 1733 0
rect 1738 -4 1742 0
rect 1748 -4 1752 0
rect 1757 -4 1761 0
rect 1773 -4 1777 0
rect 1782 -4 1786 0
rect 1792 -4 1796 0
rect 1801 -4 1805 0
rect 2091 60 2095 64
rect 2100 60 2104 64
rect 2110 60 2114 64
rect 2119 60 2123 64
rect 2135 60 2139 64
rect 2144 60 2148 64
rect 2154 60 2158 64
rect 2163 60 2167 64
rect 2228 56 2232 60
rect 2237 56 2241 60
rect 2247 56 2251 60
rect 2256 56 2260 60
rect 2272 56 2276 60
rect 2281 56 2285 60
rect 2291 56 2295 60
rect 2300 56 2304 60
rect 1880 -5 1884 -1
rect 1889 -5 1893 -1
rect 1899 -5 1903 -1
rect 1908 -5 1912 -1
rect 1924 -5 1928 -1
rect 1933 -5 1937 -1
rect 1943 -5 1947 -1
rect 1952 -5 1956 -1
rect 2166 -4 2170 0
rect 2174 -4 2178 0
rect 2121 -8 2125 -4
rect 2147 -11 2151 -7
rect 2386 5 2390 9
rect 2394 5 2398 9
rect 2343 -9 2347 -5
rect 2355 -4 2359 0
rect 2366 -9 2370 -5
rect 2268 -14 2272 -10
rect 2276 -14 2280 -10
rect 2223 -18 2227 -14
rect 2249 -21 2253 -17
rect 105 -123 109 -119
rect 113 -123 117 -119
rect 426 -146 430 -142
rect 434 -146 438 -142
rect 372 -150 376 -146
rect 383 -150 387 -146
rect 398 -150 402 -146
rect 409 -153 413 -149
rect 1245 -84 1249 -80
rect 1253 -84 1257 -80
rect 1200 -88 1204 -84
rect 1226 -91 1230 -87
rect 580 -168 584 -164
rect 588 -168 592 -164
rect 730 -168 734 -164
rect 738 -168 742 -164
rect 868 -168 872 -164
rect 876 -168 880 -164
rect 1014 -168 1018 -164
rect 1022 -168 1026 -164
rect 1138 -168 1142 -164
rect 1146 -168 1150 -164
rect 1363 -168 1367 -164
rect 1371 -168 1375 -164
rect 1510 -168 1514 -164
rect 1518 -168 1522 -164
rect 1649 -168 1653 -164
rect 1657 -168 1661 -164
rect 1773 -168 1777 -164
rect 1781 -168 1785 -164
rect 685 -172 689 -168
rect 105 -178 109 -174
rect 113 -178 117 -174
rect 537 -182 541 -178
rect 549 -177 553 -173
rect 711 -175 715 -171
rect 823 -172 827 -168
rect 849 -175 853 -171
rect 969 -172 973 -168
rect 995 -175 999 -171
rect 1093 -172 1097 -168
rect 1119 -175 1123 -171
rect 1318 -172 1322 -168
rect 1344 -175 1348 -171
rect 1465 -172 1469 -168
rect 1491 -175 1495 -171
rect 1604 -172 1608 -168
rect 1630 -175 1634 -171
rect 1728 -172 1732 -168
rect 1754 -175 1758 -171
rect 560 -182 564 -178
rect 426 -215 430 -211
rect 434 -215 438 -211
rect 372 -219 376 -215
rect 383 -219 387 -215
rect 398 -219 402 -215
rect 409 -222 413 -218
rect 3210 495 3214 499
rect 3285 495 3289 499
rect 3295 495 3299 499
rect 3311 501 3315 505
rect 426 -281 430 -277
rect 434 -281 438 -277
rect 372 -285 376 -281
rect 383 -285 387 -281
rect 398 -285 402 -281
rect 409 -288 413 -284
rect 725 -301 729 -297
rect 733 -301 737 -297
rect 680 -305 684 -301
rect 706 -308 710 -304
rect 426 -347 430 -343
rect 434 -347 438 -343
rect 372 -351 376 -347
rect 383 -351 387 -347
rect 398 -351 402 -347
rect 409 -354 413 -350
rect 863 -301 867 -297
rect 871 -301 875 -297
rect 818 -305 822 -301
rect 844 -308 848 -304
rect 1009 -301 1013 -297
rect 1017 -301 1021 -297
rect 964 -305 968 -301
rect 990 -308 994 -304
rect 1133 -301 1137 -297
rect 1141 -301 1145 -297
rect 1088 -305 1092 -301
rect 1114 -308 1118 -304
rect 1358 -301 1362 -297
rect 1366 -301 1370 -297
rect 1313 -305 1317 -301
rect 1339 -308 1343 -304
rect 1505 -301 1509 -297
rect 1513 -301 1517 -297
rect 1460 -305 1464 -301
rect 1486 -308 1490 -304
rect 1644 -301 1648 -297
rect 1652 -301 1656 -297
rect 1599 -305 1603 -301
rect 1625 -308 1629 -304
rect 1768 -301 1772 -297
rect 1776 -301 1780 -297
rect 1723 -305 1727 -301
rect 1749 -308 1753 -304
rect 721 -440 725 -436
rect 729 -440 733 -436
rect 676 -444 680 -440
rect 702 -447 706 -443
rect 859 -440 863 -436
rect 867 -440 871 -436
rect 1005 -440 1009 -436
rect 1013 -440 1017 -436
rect 1129 -440 1133 -436
rect 1137 -440 1141 -436
rect 1354 -440 1358 -436
rect 1362 -440 1366 -436
rect 814 -444 818 -440
rect 840 -447 844 -443
rect 960 -444 964 -440
rect 986 -447 990 -443
rect 1084 -444 1088 -440
rect 1110 -447 1114 -443
rect 1309 -444 1313 -440
rect 1335 -447 1339 -443
rect 1501 -440 1505 -436
rect 1509 -440 1513 -436
rect 1456 -444 1460 -440
rect 1482 -447 1486 -443
rect 1640 -440 1644 -436
rect 1648 -440 1652 -436
rect 1595 -444 1599 -440
rect 1621 -447 1625 -443
rect 1764 -440 1768 -436
rect 1772 -440 1776 -436
rect 1719 -444 1723 -440
rect 1745 -447 1749 -443
rect 1880 -484 1884 -480
rect 1888 -484 1892 -480
rect 1835 -488 1839 -484
rect 1861 -491 1865 -487
rect 2968 452 2972 456
rect 2976 452 2980 456
rect 3660 450 3664 454
rect 3673 453 3677 457
rect 3686 450 3690 454
rect 3699 453 3703 457
rect 3712 453 3716 457
rect 3720 453 3724 457
rect 3733 453 3737 457
rect 3341 395 3345 399
rect 3403 395 3407 399
rect 3412 395 3416 399
rect 3428 401 3432 405
rect 2970 386 2974 390
rect 2978 386 2982 390
rect 2973 319 2977 323
rect 2981 319 2985 323
rect 2973 252 2977 256
rect 2981 252 2985 256
rect 2991 147 2995 151
rect 2999 147 3003 151
rect 2891 103 2895 107
rect 2900 103 2904 107
rect 2910 103 2914 107
rect 2919 103 2923 107
rect 2935 103 2939 107
rect 2944 103 2948 107
rect 2954 103 2958 107
rect 2963 103 2967 107
rect 2993 -14 2997 -10
rect 3001 -14 3005 -10
rect 2893 -58 2897 -54
rect 2902 -58 2906 -54
rect 2912 -58 2916 -54
rect 2921 -58 2925 -54
rect 2937 -58 2941 -54
rect 2946 -58 2950 -54
rect 2956 -58 2960 -54
rect 2965 -58 2969 -54
rect 3479 357 3483 361
rect 3529 357 3533 361
rect 3538 357 3542 361
rect 3554 363 3558 367
rect 3656 329 3660 333
rect 3664 329 3668 333
rect 3608 325 3612 329
rect 3640 322 3644 326
rect 3762 -69 3766 -65
rect 3770 -69 3774 -65
rect 3588 -79 3592 -75
rect 3650 -79 3654 -75
rect 3659 -79 3663 -75
rect 3675 -73 3679 -69
rect 3703 -73 3707 -69
rect 3740 -76 3744 -72
rect 2992 -168 2996 -164
rect 3000 -168 3004 -164
rect 2892 -212 2896 -208
rect 2901 -212 2905 -208
rect 2911 -212 2915 -208
rect 2920 -212 2924 -208
rect 2936 -212 2940 -208
rect 2945 -212 2949 -208
rect 2955 -212 2959 -208
rect 2964 -212 2968 -208
rect 2992 -316 2996 -312
rect 3000 -316 3004 -312
rect 3651 -330 3655 -326
rect 3664 -327 3668 -323
rect 3677 -330 3681 -326
rect 3690 -327 3694 -323
rect 3703 -327 3707 -323
rect 3711 -327 3715 -323
rect 3724 -327 3728 -323
rect 2892 -360 2896 -356
rect 2901 -360 2905 -356
rect 2911 -360 2915 -356
rect 2920 -360 2924 -356
rect 2936 -360 2940 -356
rect 2945 -360 2949 -356
rect 2955 -360 2959 -356
rect 2964 -360 2968 -356
rect 3425 -394 3429 -390
rect 3500 -394 3504 -390
rect 3510 -394 3514 -390
rect 3526 -388 3530 -384
rect 2968 -443 2972 -439
rect 2976 -443 2980 -439
rect 3293 -478 3297 -474
rect 3355 -478 3359 -474
rect 3364 -478 3368 -474
rect 3380 -472 3384 -468
rect 2970 -509 2974 -505
rect 2978 -509 2982 -505
rect 3152 -553 3156 -549
rect 3202 -553 3206 -549
rect 3211 -553 3215 -549
rect 3227 -547 3231 -543
rect 2973 -576 2977 -572
rect 2981 -576 2985 -572
rect 1880 -589 1884 -585
rect 1888 -589 1892 -585
rect 1835 -593 1839 -589
rect 1861 -596 1865 -592
rect 3105 -615 3109 -611
rect 3113 -615 3117 -611
rect 3057 -619 3061 -615
rect 3089 -622 3093 -618
rect 2973 -643 2977 -639
rect 2981 -643 2985 -639
rect 1880 -711 1884 -707
rect 1888 -711 1892 -707
rect 1835 -715 1839 -711
rect 1861 -718 1865 -714
rect 1880 -818 1884 -814
rect 1888 -818 1892 -814
rect 1835 -822 1839 -818
rect 1861 -825 1865 -821
<< pdcontact >>
rect 2093 931 2097 935
rect 2102 931 2106 935
rect 2112 931 2116 935
rect 2121 931 2125 935
rect 2137 931 2141 935
rect 2146 931 2150 935
rect 2156 931 2160 935
rect 2165 931 2169 935
rect 2230 927 2234 931
rect 2239 927 2243 931
rect 2249 927 2253 931
rect 2258 927 2262 931
rect 2274 927 2278 931
rect 2283 927 2287 931
rect 2293 927 2297 931
rect 2302 927 2306 931
rect 2345 869 2349 873
rect 2388 869 2392 873
rect 2396 869 2400 873
rect 2368 864 2372 868
rect 2123 859 2127 863
rect 2135 860 2139 864
rect 2149 859 2153 863
rect 2168 860 2172 864
rect 2176 860 2180 864
rect 2225 849 2229 853
rect 2237 850 2241 854
rect 2251 849 2255 853
rect 2270 850 2274 854
rect 2278 850 2282 854
rect 2091 655 2095 659
rect 2100 655 2104 659
rect 2110 655 2114 659
rect 2119 655 2123 659
rect 2135 655 2139 659
rect 2144 655 2148 659
rect 2154 655 2158 659
rect 2163 655 2167 659
rect 2228 651 2232 655
rect 2237 651 2241 655
rect 2247 651 2251 655
rect 2256 651 2260 655
rect 2272 651 2276 655
rect 2281 651 2285 655
rect 2291 651 2295 655
rect 2300 651 2304 655
rect 2343 593 2347 597
rect 2386 593 2390 597
rect 2394 593 2398 597
rect 2366 588 2370 592
rect 2121 583 2125 587
rect 2133 584 2137 588
rect 2147 583 2151 587
rect 2166 584 2170 588
rect 2174 584 2178 588
rect 2223 573 2227 577
rect 2235 574 2239 578
rect 2249 573 2253 577
rect 2268 574 2272 578
rect 2276 574 2280 578
rect 2088 376 2092 380
rect 2097 376 2101 380
rect 2107 376 2111 380
rect 2116 376 2120 380
rect 2132 376 2136 380
rect 2141 376 2145 380
rect 2151 376 2155 380
rect 2160 376 2164 380
rect 2225 372 2229 376
rect 2234 372 2238 376
rect 2244 372 2248 376
rect 2253 372 2257 376
rect 2269 372 2273 376
rect 2278 372 2282 376
rect 2288 372 2292 376
rect 2297 372 2301 376
rect 2340 314 2344 318
rect 2383 314 2387 318
rect 2391 314 2395 318
rect 2363 309 2367 313
rect 2118 304 2122 308
rect 2130 305 2134 309
rect 2144 304 2148 308
rect 2163 305 2167 309
rect 2171 305 2175 309
rect 2220 294 2224 298
rect 2232 295 2236 299
rect 2246 294 2250 298
rect 2265 295 2269 299
rect 2273 295 2277 299
rect 1428 30 1432 34
rect 1437 30 1441 34
rect 1447 30 1451 34
rect 1456 30 1460 34
rect 1472 30 1476 34
rect 1481 30 1485 34
rect 1491 30 1495 34
rect 1500 30 1504 34
rect 1577 28 1581 32
rect 1586 28 1590 32
rect 1596 28 1600 32
rect 1605 28 1609 32
rect 1621 28 1625 32
rect 1630 28 1634 32
rect 1640 28 1644 32
rect 1649 28 1653 32
rect 1729 27 1733 31
rect 1738 27 1742 31
rect 1748 27 1752 31
rect 1757 27 1761 31
rect 1773 27 1777 31
rect 1782 27 1786 31
rect 1792 27 1796 31
rect 1801 27 1805 31
rect 2091 91 2095 95
rect 2100 91 2104 95
rect 2110 91 2114 95
rect 2119 91 2123 95
rect 2135 91 2139 95
rect 2144 91 2148 95
rect 2154 91 2158 95
rect 2163 91 2167 95
rect 2228 87 2232 91
rect 2237 87 2241 91
rect 2247 87 2251 91
rect 2256 87 2260 91
rect 2272 87 2276 91
rect 2281 87 2285 91
rect 2291 87 2295 91
rect 2300 87 2304 91
rect 1880 26 1884 30
rect 1889 26 1893 30
rect 1899 26 1903 30
rect 1908 26 1912 30
rect 1924 26 1928 30
rect 1933 26 1937 30
rect 1943 26 1947 30
rect 1952 26 1956 30
rect 2343 29 2347 33
rect 2386 29 2390 33
rect 2394 29 2398 33
rect 2366 24 2370 28
rect 2121 19 2125 23
rect 2133 20 2137 24
rect 2147 19 2151 23
rect 2166 20 2170 24
rect 2174 20 2178 24
rect 2223 9 2227 13
rect 2235 10 2239 14
rect 2249 9 2253 13
rect 2268 10 2272 14
rect 2276 10 2280 14
rect 1200 -61 1204 -57
rect 1212 -60 1216 -56
rect 1226 -61 1230 -57
rect 1245 -60 1249 -56
rect 1253 -60 1257 -56
rect 105 -99 109 -95
rect 113 -99 117 -95
rect 372 -123 376 -119
rect 383 -122 387 -118
rect 398 -123 402 -119
rect 409 -122 413 -118
rect 426 -122 430 -118
rect 434 -122 438 -118
rect 105 -154 109 -150
rect 113 -154 117 -150
rect 537 -144 541 -140
rect 580 -144 584 -140
rect 588 -144 592 -140
rect 560 -149 564 -145
rect 685 -145 689 -141
rect 697 -144 701 -140
rect 711 -145 715 -141
rect 730 -144 734 -140
rect 738 -144 742 -140
rect 823 -145 827 -141
rect 835 -144 839 -140
rect 849 -145 853 -141
rect 868 -144 872 -140
rect 876 -144 880 -140
rect 969 -145 973 -141
rect 981 -144 985 -140
rect 995 -145 999 -141
rect 1014 -144 1018 -140
rect 1022 -144 1026 -140
rect 1093 -145 1097 -141
rect 1105 -144 1109 -140
rect 1119 -145 1123 -141
rect 1138 -144 1142 -140
rect 1146 -144 1150 -140
rect 1318 -145 1322 -141
rect 1330 -144 1334 -140
rect 1344 -145 1348 -141
rect 1363 -144 1367 -140
rect 1371 -144 1375 -140
rect 1465 -145 1469 -141
rect 1477 -144 1481 -140
rect 1491 -145 1495 -141
rect 1510 -144 1514 -140
rect 1518 -144 1522 -140
rect 1604 -145 1608 -141
rect 1616 -144 1620 -140
rect 1630 -145 1634 -141
rect 1649 -144 1653 -140
rect 1657 -144 1661 -140
rect 1728 -145 1732 -141
rect 1740 -144 1744 -140
rect 1754 -145 1758 -141
rect 1773 -144 1777 -140
rect 1781 -144 1785 -140
rect 372 -192 376 -188
rect 383 -191 387 -187
rect 398 -192 402 -188
rect 409 -191 413 -187
rect 426 -191 430 -187
rect 434 -191 438 -187
rect 372 -258 376 -254
rect 383 -257 387 -253
rect 398 -258 402 -254
rect 409 -257 413 -253
rect 426 -257 430 -253
rect 434 -257 438 -253
rect 3210 530 3214 534
rect 3223 530 3227 534
rect 3240 530 3244 534
rect 3255 530 3259 534
rect 3270 530 3274 534
rect 3285 530 3289 534
rect 3295 530 3299 534
rect 3311 530 3315 534
rect 2968 476 2972 480
rect 2976 476 2980 480
rect 680 -278 684 -274
rect 692 -277 696 -273
rect 706 -278 710 -274
rect 725 -277 729 -273
rect 733 -277 737 -273
rect 818 -278 822 -274
rect 830 -277 834 -273
rect 844 -278 848 -274
rect 863 -277 867 -273
rect 871 -277 875 -273
rect 372 -324 376 -320
rect 383 -323 387 -319
rect 398 -324 402 -320
rect 409 -323 413 -319
rect 426 -323 430 -319
rect 434 -323 438 -319
rect 964 -278 968 -274
rect 976 -277 980 -273
rect 990 -278 994 -274
rect 1009 -277 1013 -273
rect 1017 -277 1021 -273
rect 1088 -278 1092 -274
rect 1100 -277 1104 -273
rect 1114 -278 1118 -274
rect 1133 -277 1137 -273
rect 1141 -277 1145 -273
rect 1313 -278 1317 -274
rect 1325 -277 1329 -273
rect 1339 -278 1343 -274
rect 1358 -277 1362 -273
rect 1366 -277 1370 -273
rect 1460 -278 1464 -274
rect 1472 -277 1476 -273
rect 1486 -278 1490 -274
rect 1505 -277 1509 -273
rect 1513 -277 1517 -273
rect 1599 -278 1603 -274
rect 1611 -277 1615 -273
rect 1625 -278 1629 -274
rect 1644 -277 1648 -273
rect 1652 -277 1656 -273
rect 1723 -278 1727 -274
rect 1735 -277 1739 -273
rect 1749 -278 1753 -274
rect 1768 -277 1772 -273
rect 1776 -277 1780 -273
rect 676 -417 680 -413
rect 688 -416 692 -412
rect 702 -417 706 -413
rect 721 -416 725 -412
rect 729 -416 733 -412
rect 814 -417 818 -413
rect 826 -416 830 -412
rect 840 -417 844 -413
rect 859 -416 863 -412
rect 867 -416 871 -412
rect 960 -417 964 -413
rect 972 -416 976 -412
rect 986 -417 990 -413
rect 1005 -416 1009 -412
rect 1013 -416 1017 -412
rect 1084 -417 1088 -413
rect 1096 -416 1100 -412
rect 1110 -417 1114 -413
rect 1129 -416 1133 -412
rect 1137 -416 1141 -412
rect 1309 -417 1313 -413
rect 1321 -416 1325 -412
rect 1335 -417 1339 -413
rect 1354 -416 1358 -412
rect 1362 -416 1366 -412
rect 1456 -417 1460 -413
rect 1468 -416 1472 -412
rect 1482 -417 1486 -413
rect 1501 -416 1505 -412
rect 1509 -416 1513 -412
rect 1595 -417 1599 -413
rect 1607 -416 1611 -412
rect 1621 -417 1625 -413
rect 1640 -416 1644 -412
rect 1648 -416 1652 -412
rect 1719 -417 1723 -413
rect 1731 -416 1735 -412
rect 1745 -417 1749 -413
rect 1764 -416 1768 -412
rect 1772 -416 1776 -412
rect 1835 -461 1839 -457
rect 1847 -460 1851 -456
rect 1861 -461 1865 -457
rect 1880 -460 1884 -456
rect 1888 -460 1892 -456
rect 1835 -566 1839 -562
rect 1847 -565 1851 -561
rect 1861 -566 1865 -562
rect 1880 -565 1884 -561
rect 1888 -565 1892 -561
rect 3341 430 3345 434
rect 3356 430 3361 434
rect 3374 430 3378 434
rect 3389 430 3393 434
rect 3403 430 3407 434
rect 3412 430 3416 434
rect 3428 430 3432 434
rect 3660 480 3664 484
rect 3712 480 3716 484
rect 3720 480 3724 484
rect 3733 480 3737 484
rect 2970 410 2974 414
rect 2978 410 2982 414
rect 2973 343 2977 347
rect 2981 343 2985 347
rect 2973 276 2977 280
rect 2981 276 2985 280
rect 2991 171 2995 175
rect 2999 171 3003 175
rect 2891 134 2895 138
rect 2900 134 2904 138
rect 2910 134 2914 138
rect 2919 134 2923 138
rect 2935 134 2939 138
rect 2944 134 2948 138
rect 2954 134 2958 138
rect 2963 134 2967 138
rect 2993 10 2997 14
rect 3001 10 3005 14
rect 2893 -27 2897 -23
rect 2902 -27 2906 -23
rect 2912 -27 2916 -23
rect 2921 -27 2925 -23
rect 2937 -27 2941 -23
rect 2946 -27 2950 -23
rect 2956 -27 2960 -23
rect 2965 -27 2969 -23
rect 3479 392 3483 396
rect 3494 392 3499 396
rect 3512 392 3516 396
rect 3529 392 3533 396
rect 3538 392 3542 396
rect 3554 392 3558 396
rect 3608 352 3612 356
rect 3619 353 3623 357
rect 3629 352 3633 356
rect 3640 353 3644 357
rect 3656 353 3660 357
rect 3664 353 3668 357
rect 3588 -44 3592 -40
rect 3603 -44 3608 -40
rect 3621 -44 3625 -40
rect 3636 -44 3640 -40
rect 3650 -44 3654 -40
rect 3659 -44 3663 -40
rect 3675 -44 3679 -40
rect 3703 -46 3707 -42
rect 3714 -45 3718 -41
rect 3729 -46 3733 -42
rect 3740 -45 3744 -41
rect 3762 -45 3766 -41
rect 3770 -45 3774 -41
rect 2992 -144 2996 -140
rect 3000 -144 3004 -140
rect 2892 -181 2896 -177
rect 2901 -181 2905 -177
rect 2911 -181 2915 -177
rect 2920 -181 2924 -177
rect 2936 -181 2940 -177
rect 2945 -181 2949 -177
rect 2955 -181 2959 -177
rect 2964 -181 2968 -177
rect 2992 -292 2996 -288
rect 3000 -292 3004 -288
rect 3651 -300 3655 -296
rect 3703 -300 3707 -296
rect 3711 -300 3715 -296
rect 3724 -300 3728 -296
rect 2892 -329 2896 -325
rect 2901 -329 2905 -325
rect 2911 -329 2915 -325
rect 2920 -329 2924 -325
rect 2936 -329 2940 -325
rect 2945 -329 2949 -325
rect 2955 -329 2959 -325
rect 2964 -329 2968 -325
rect 3425 -359 3429 -355
rect 3438 -359 3442 -355
rect 3455 -359 3459 -355
rect 3470 -359 3474 -355
rect 3485 -359 3489 -355
rect 3500 -359 3504 -355
rect 3510 -359 3514 -355
rect 3526 -359 3530 -355
rect 2968 -419 2972 -415
rect 2976 -419 2980 -415
rect 3293 -443 3297 -439
rect 3308 -443 3313 -439
rect 3326 -443 3330 -439
rect 3341 -443 3345 -439
rect 3355 -443 3359 -439
rect 3364 -443 3368 -439
rect 3380 -443 3384 -439
rect 2970 -485 2974 -481
rect 2978 -485 2982 -481
rect 3152 -518 3156 -514
rect 3167 -518 3172 -514
rect 3185 -518 3189 -514
rect 3202 -518 3206 -514
rect 3211 -518 3215 -514
rect 3227 -518 3231 -514
rect 2973 -552 2977 -548
rect 2981 -552 2985 -548
rect 3057 -592 3061 -588
rect 3068 -591 3072 -587
rect 3078 -592 3082 -588
rect 3089 -591 3093 -587
rect 3105 -591 3109 -587
rect 3113 -591 3117 -587
rect 2973 -619 2977 -615
rect 2981 -619 2985 -615
rect 1835 -688 1839 -684
rect 1847 -687 1851 -683
rect 1861 -688 1865 -684
rect 1880 -687 1884 -683
rect 1888 -687 1892 -683
rect 1835 -795 1839 -791
rect 1847 -794 1851 -790
rect 1861 -795 1865 -791
rect 1880 -794 1884 -790
rect 1888 -794 1892 -790
<< polysilicon >>
rect 2083 965 2119 967
rect 2083 880 2085 965
rect 2098 936 2100 939
rect 2117 936 2119 965
rect 2220 961 2256 963
rect 2142 936 2144 939
rect 2161 936 2163 939
rect 2098 919 2100 931
rect 2117 928 2119 931
rect 2142 919 2144 931
rect 2098 917 2119 919
rect 2098 905 2100 908
rect 2117 905 2119 917
rect 2143 915 2144 919
rect 2142 905 2144 915
rect 2161 905 2163 931
rect 2172 916 2178 918
rect 2098 880 2100 900
rect 2117 889 2119 900
rect 2142 897 2144 900
rect 2161 889 2163 900
rect 2121 887 2163 889
rect 2176 880 2178 916
rect 2083 878 2178 880
rect 2220 875 2222 961
rect 2235 932 2237 935
rect 2254 932 2256 961
rect 2279 932 2281 935
rect 2298 932 2300 935
rect 2235 915 2237 927
rect 2254 924 2256 927
rect 2279 915 2281 927
rect 2235 913 2256 915
rect 2235 901 2237 904
rect 2254 901 2256 913
rect 2280 911 2281 915
rect 2279 901 2281 911
rect 2298 901 2300 927
rect 2309 912 2315 914
rect 2235 875 2237 896
rect 2254 886 2256 896
rect 2279 893 2281 896
rect 2298 885 2300 896
rect 2256 883 2300 885
rect 2313 875 2315 912
rect 2220 873 2315 875
rect 2353 873 2355 876
rect 2362 873 2364 876
rect 2393 873 2395 876
rect 2129 864 2131 867
rect 2144 864 2146 867
rect 2173 864 2175 867
rect 2129 852 2131 859
rect 2129 836 2131 848
rect 2144 843 2146 859
rect 2173 847 2175 860
rect 2353 858 2355 864
rect 2231 854 2233 857
rect 2246 854 2248 857
rect 2275 854 2277 857
rect 2344 855 2355 858
rect 2168 845 2175 847
rect 2134 840 2135 843
rect 2139 840 2146 843
rect 2173 840 2175 845
rect 2231 842 2233 849
rect 2144 836 2146 840
rect 2173 833 2175 836
rect 2129 826 2131 829
rect 2144 826 2146 829
rect 2213 806 2215 838
rect 2231 826 2233 838
rect 2246 833 2248 849
rect 2275 837 2277 850
rect 2353 840 2355 855
rect 2362 851 2364 864
rect 2393 856 2395 869
rect 2388 854 2395 856
rect 2363 847 2364 851
rect 2393 849 2395 854
rect 2405 853 2442 857
rect 2362 840 2364 847
rect 2393 842 2395 845
rect 2270 835 2277 837
rect 2236 830 2237 833
rect 2241 830 2248 833
rect 2275 830 2277 835
rect 2246 826 2248 830
rect 2353 828 2355 831
rect 2362 828 2364 831
rect 2275 823 2277 826
rect 2231 816 2233 819
rect 2246 816 2248 819
rect 2081 689 2117 691
rect 2081 604 2083 689
rect 2096 660 2098 663
rect 2115 660 2117 689
rect 2218 685 2254 687
rect 2140 660 2142 663
rect 2159 660 2161 663
rect 2096 643 2098 655
rect 2115 652 2117 655
rect 2140 643 2142 655
rect 2096 641 2117 643
rect 2096 629 2098 632
rect 2115 629 2117 641
rect 2141 639 2142 643
rect 2140 629 2142 639
rect 2159 629 2161 655
rect 2170 640 2176 642
rect 2096 604 2098 624
rect 2115 613 2117 624
rect 2140 621 2142 624
rect 2159 613 2161 624
rect 2119 611 2161 613
rect 2174 604 2176 640
rect 2081 602 2176 604
rect 2218 599 2220 685
rect 2233 656 2235 659
rect 2252 656 2254 685
rect 2277 656 2279 659
rect 2296 656 2298 659
rect 2233 639 2235 651
rect 2252 648 2254 651
rect 2277 639 2279 651
rect 2233 637 2254 639
rect 2233 625 2235 628
rect 2252 625 2254 637
rect 2278 635 2279 639
rect 2277 625 2279 635
rect 2296 625 2298 651
rect 2307 636 2313 638
rect 2233 599 2235 620
rect 2252 610 2254 620
rect 2277 617 2279 620
rect 2296 609 2298 620
rect 2254 607 2298 609
rect 2311 599 2313 636
rect 2218 597 2313 599
rect 2351 597 2353 600
rect 2360 597 2362 600
rect 2391 597 2393 600
rect 2127 588 2129 591
rect 2142 588 2144 591
rect 2171 588 2173 591
rect 2127 576 2129 583
rect 2127 560 2129 572
rect 2142 567 2144 583
rect 2171 571 2173 584
rect 2351 582 2353 588
rect 2229 578 2231 581
rect 2244 578 2246 581
rect 2273 578 2275 581
rect 2342 579 2353 582
rect 2166 569 2173 571
rect 2132 564 2133 567
rect 2137 564 2144 567
rect 2171 564 2173 569
rect 2229 566 2231 573
rect 2142 560 2144 564
rect 2171 557 2173 560
rect 2127 550 2129 553
rect 2142 550 2144 553
rect 2211 516 2213 562
rect 2229 550 2231 562
rect 2244 557 2246 573
rect 2273 561 2275 574
rect 2351 564 2353 579
rect 2360 575 2362 588
rect 2391 580 2393 593
rect 2386 578 2393 580
rect 2361 571 2362 575
rect 2391 573 2393 578
rect 2360 564 2362 571
rect 2391 566 2393 569
rect 2268 559 2275 561
rect 2234 554 2235 557
rect 2239 554 2246 557
rect 2273 554 2275 559
rect 2244 550 2246 554
rect 2351 552 2353 555
rect 2360 552 2362 555
rect 2273 547 2275 550
rect 2229 540 2231 543
rect 2244 540 2246 543
rect 2439 516 2442 853
rect 2211 513 2442 516
rect 2748 575 3759 577
rect 2078 410 2114 412
rect 2078 325 2080 410
rect 2093 381 2095 384
rect 2112 381 2114 410
rect 2215 406 2251 408
rect 2137 381 2139 384
rect 2156 381 2158 384
rect 2093 364 2095 376
rect 2112 373 2114 376
rect 2137 364 2139 376
rect 2093 362 2114 364
rect 2093 350 2095 353
rect 2112 350 2114 362
rect 2138 360 2139 364
rect 2137 350 2139 360
rect 2156 350 2158 376
rect 2167 361 2173 363
rect 2093 325 2095 345
rect 2112 334 2114 345
rect 2137 342 2139 345
rect 2156 334 2158 345
rect 2116 332 2158 334
rect 2171 325 2173 361
rect 2078 323 2173 325
rect 2215 320 2217 406
rect 2230 377 2232 380
rect 2249 377 2251 406
rect 2274 377 2276 380
rect 2293 377 2295 380
rect 2230 360 2232 372
rect 2249 369 2251 372
rect 2274 360 2276 372
rect 2230 358 2251 360
rect 2230 346 2232 349
rect 2249 346 2251 358
rect 2275 356 2276 360
rect 2274 346 2276 356
rect 2293 346 2295 372
rect 2304 357 2310 359
rect 2230 320 2232 341
rect 2249 331 2251 341
rect 2274 338 2276 341
rect 2293 330 2295 341
rect 2251 328 2295 330
rect 2308 320 2310 357
rect 2215 318 2310 320
rect 2348 318 2350 321
rect 2357 318 2359 321
rect 2388 318 2390 321
rect 2124 309 2126 312
rect 2139 309 2141 312
rect 2168 309 2170 312
rect 2124 297 2126 304
rect 2124 281 2126 293
rect 2139 288 2141 304
rect 2168 292 2170 305
rect 2348 303 2350 309
rect 2226 299 2228 302
rect 2241 299 2243 302
rect 2270 299 2272 302
rect 2339 300 2350 303
rect 2163 290 2170 292
rect 2129 285 2130 288
rect 2134 285 2141 288
rect 2168 285 2170 290
rect 2226 287 2228 294
rect 2139 281 2141 285
rect 2168 278 2170 281
rect 2124 271 2126 274
rect 2139 271 2141 274
rect 2208 251 2210 283
rect 2226 271 2228 283
rect 2241 278 2243 294
rect 2270 282 2272 295
rect 2348 285 2350 300
rect 2357 296 2359 309
rect 2388 301 2390 314
rect 2383 299 2390 301
rect 2358 292 2359 296
rect 2388 294 2390 299
rect 2400 298 2430 302
rect 2357 285 2359 292
rect 2388 287 2390 290
rect 2265 280 2272 282
rect 2231 275 2232 278
rect 2236 275 2243 278
rect 2270 275 2272 280
rect 2241 271 2243 275
rect 2348 273 2350 276
rect 2357 273 2359 276
rect 2270 268 2272 271
rect 2226 261 2228 264
rect 2241 261 2243 264
rect 2081 125 2117 127
rect 1418 64 1454 66
rect 1418 -21 1420 64
rect 1433 35 1435 38
rect 1452 35 1454 64
rect 1567 62 1603 64
rect 1477 35 1479 38
rect 1496 35 1498 38
rect 1433 18 1435 30
rect 1452 27 1454 30
rect 1477 18 1479 30
rect 1433 16 1454 18
rect 1433 4 1435 7
rect 1452 4 1454 16
rect 1478 14 1479 18
rect 1477 4 1479 14
rect 1496 4 1498 30
rect 1507 15 1513 17
rect 1433 -21 1435 -1
rect 1452 -12 1454 -1
rect 1477 -4 1479 -1
rect 1496 -12 1498 -1
rect 1456 -14 1498 -12
rect 1511 -21 1513 15
rect 1418 -23 1513 -21
rect 1567 -23 1569 62
rect 1582 33 1584 36
rect 1601 33 1603 62
rect 1719 61 1755 63
rect 1626 33 1628 36
rect 1645 33 1647 36
rect 1582 16 1584 28
rect 1601 25 1603 28
rect 1626 16 1628 28
rect 1582 14 1603 16
rect 1582 2 1584 5
rect 1601 2 1603 14
rect 1627 12 1628 16
rect 1626 2 1628 12
rect 1645 2 1647 28
rect 1656 13 1662 15
rect 1582 -23 1584 -3
rect 1601 -14 1603 -3
rect 1626 -6 1628 -3
rect 1645 -14 1647 -3
rect 1605 -16 1647 -14
rect 1660 -23 1662 13
rect 1567 -25 1662 -23
rect 1719 -24 1721 61
rect 1734 32 1736 35
rect 1753 32 1755 61
rect 1870 60 1906 62
rect 1778 32 1780 35
rect 1797 32 1799 35
rect 1734 15 1736 27
rect 1753 24 1755 27
rect 1778 15 1780 27
rect 1734 13 1755 15
rect 1734 1 1736 4
rect 1753 1 1755 13
rect 1779 11 1780 15
rect 1778 1 1780 11
rect 1797 1 1799 27
rect 1808 12 1814 14
rect 1734 -24 1736 -4
rect 1753 -15 1755 -4
rect 1778 -7 1780 -4
rect 1797 -15 1799 -4
rect 1757 -17 1799 -15
rect 1812 -24 1814 12
rect 1719 -26 1814 -24
rect 1870 -25 1872 60
rect 1885 31 1887 34
rect 1904 31 1906 60
rect 2081 40 2083 125
rect 2096 96 2098 99
rect 2115 96 2117 125
rect 2218 121 2254 123
rect 2140 96 2142 99
rect 2159 96 2161 99
rect 2096 79 2098 91
rect 2115 88 2117 91
rect 2140 79 2142 91
rect 2096 77 2117 79
rect 2096 65 2098 68
rect 2115 65 2117 77
rect 2141 75 2142 79
rect 2140 65 2142 75
rect 2159 65 2161 91
rect 2170 76 2176 78
rect 2096 40 2098 60
rect 2115 49 2117 60
rect 2140 57 2142 60
rect 2159 49 2161 60
rect 2119 47 2161 49
rect 2174 40 2176 76
rect 2081 38 2176 40
rect 2218 35 2220 121
rect 2233 92 2235 95
rect 2252 92 2254 121
rect 2277 92 2279 95
rect 2296 92 2298 95
rect 2233 75 2235 87
rect 2252 84 2254 87
rect 2277 75 2279 87
rect 2233 73 2254 75
rect 2233 61 2235 64
rect 2252 61 2254 73
rect 2278 71 2279 75
rect 2277 61 2279 71
rect 2296 61 2298 87
rect 2307 72 2313 74
rect 2233 35 2235 56
rect 2252 46 2254 56
rect 2277 53 2279 56
rect 2296 45 2298 56
rect 2254 43 2298 45
rect 2311 35 2313 72
rect 1929 31 1931 34
rect 1948 31 1950 34
rect 2218 33 2313 35
rect 2351 33 2353 36
rect 2360 33 2362 36
rect 2391 33 2393 36
rect 1885 14 1887 26
rect 1904 23 1906 26
rect 1929 14 1931 26
rect 1885 12 1906 14
rect 1885 0 1887 3
rect 1904 0 1906 12
rect 1930 10 1931 14
rect 1929 0 1931 10
rect 1948 0 1950 26
rect 2127 24 2129 27
rect 2142 24 2144 27
rect 2171 24 2173 27
rect 1959 11 1965 13
rect 2127 12 2129 19
rect 1885 -25 1887 -5
rect 1904 -16 1906 -5
rect 1929 -8 1931 -5
rect 1948 -16 1950 -5
rect 1908 -18 1950 -16
rect 1963 -25 1965 11
rect 2127 -4 2129 8
rect 2142 3 2144 19
rect 2171 7 2173 20
rect 2351 18 2353 24
rect 2229 14 2231 17
rect 2244 14 2246 17
rect 2273 14 2275 17
rect 2342 15 2353 18
rect 2166 5 2173 7
rect 2132 0 2133 3
rect 2137 0 2144 3
rect 2171 0 2173 5
rect 2229 2 2231 9
rect 2142 -4 2144 0
rect 2171 -7 2173 -4
rect 2127 -14 2129 -11
rect 2142 -14 2144 -11
rect 1870 -27 1965 -25
rect 2211 -36 2213 -2
rect 2229 -14 2231 -2
rect 2244 -7 2246 9
rect 2273 -3 2275 10
rect 2351 0 2353 15
rect 2360 11 2362 24
rect 2391 16 2393 29
rect 2386 14 2393 16
rect 2361 7 2362 11
rect 2391 9 2393 14
rect 2360 0 2362 7
rect 2391 2 2393 5
rect 2268 -5 2275 -3
rect 2234 -10 2235 -7
rect 2239 -10 2246 -7
rect 2273 -10 2275 -5
rect 2244 -14 2246 -10
rect 2351 -12 2353 -9
rect 2360 -12 2362 -9
rect 2273 -17 2275 -14
rect 2229 -24 2231 -21
rect 2244 -24 2246 -21
rect 2428 -36 2430 298
rect 2211 -38 2430 -36
rect 1206 -56 1208 -53
rect 1221 -56 1223 -53
rect 1250 -56 1252 -53
rect 1206 -68 1208 -61
rect 1171 -72 1208 -68
rect 1171 -77 1173 -72
rect 518 -79 1173 -77
rect 110 -95 112 -92
rect 110 -112 112 -99
rect 105 -114 112 -112
rect 110 -119 112 -114
rect 378 -118 380 -115
rect 404 -118 406 -115
rect 431 -118 433 -115
rect 110 -126 112 -123
rect 378 -132 380 -123
rect 404 -132 406 -123
rect 378 -146 380 -136
rect 404 -146 406 -136
rect 431 -135 433 -122
rect 426 -137 433 -135
rect 431 -142 433 -137
rect 110 -150 112 -147
rect 431 -149 433 -146
rect 110 -167 112 -154
rect 378 -156 380 -153
rect 404 -156 406 -153
rect 518 -163 520 -79
rect 1195 -81 1198 -77
rect 1195 -125 1197 -81
rect 1206 -84 1208 -72
rect 1221 -77 1223 -61
rect 1250 -73 1252 -60
rect 1245 -75 1252 -73
rect 1211 -80 1212 -77
rect 1216 -80 1223 -77
rect 1250 -80 1252 -75
rect 1221 -84 1223 -80
rect 1250 -87 1252 -84
rect 1206 -94 1208 -91
rect 1221 -94 1223 -91
rect 601 -127 1720 -125
rect 545 -140 547 -137
rect 554 -140 556 -137
rect 585 -140 587 -137
rect 545 -155 547 -149
rect 536 -158 547 -155
rect 105 -169 112 -167
rect 110 -174 112 -169
rect 545 -173 547 -158
rect 554 -162 556 -149
rect 585 -157 587 -144
rect 601 -156 604 -127
rect 674 -152 676 -127
rect 691 -140 693 -137
rect 706 -140 708 -137
rect 735 -140 737 -137
rect 691 -152 693 -145
rect 674 -156 693 -152
rect 580 -159 587 -157
rect 555 -166 556 -162
rect 585 -164 587 -159
rect 597 -160 604 -156
rect 554 -173 556 -166
rect 691 -168 693 -156
rect 706 -161 708 -145
rect 735 -157 737 -144
rect 812 -152 814 -127
rect 829 -140 831 -137
rect 844 -140 846 -137
rect 873 -140 875 -137
rect 829 -152 831 -145
rect 812 -156 831 -152
rect 730 -159 737 -157
rect 696 -164 697 -161
rect 701 -164 708 -161
rect 735 -164 737 -159
rect 706 -168 708 -164
rect 829 -168 831 -156
rect 844 -161 846 -145
rect 873 -157 875 -144
rect 958 -152 960 -127
rect 975 -140 977 -137
rect 990 -140 992 -137
rect 1019 -140 1021 -137
rect 975 -152 977 -145
rect 958 -156 977 -152
rect 868 -159 875 -157
rect 834 -164 835 -161
rect 839 -164 846 -161
rect 873 -164 875 -159
rect 844 -168 846 -164
rect 975 -168 977 -156
rect 990 -161 992 -145
rect 1019 -157 1021 -144
rect 1082 -152 1084 -127
rect 1099 -140 1101 -137
rect 1114 -140 1116 -137
rect 1143 -140 1145 -137
rect 1099 -152 1101 -145
rect 1082 -156 1101 -152
rect 1014 -159 1021 -157
rect 980 -164 981 -161
rect 985 -164 992 -161
rect 1019 -164 1021 -159
rect 990 -168 992 -164
rect 1099 -168 1101 -156
rect 1114 -161 1116 -145
rect 1143 -157 1145 -144
rect 1306 -152 1308 -127
rect 1324 -140 1326 -137
rect 1339 -140 1341 -137
rect 1368 -140 1370 -137
rect 1324 -152 1326 -145
rect 1306 -156 1326 -152
rect 1138 -159 1145 -157
rect 1104 -164 1105 -161
rect 1109 -164 1116 -161
rect 1143 -164 1145 -159
rect 1114 -168 1116 -164
rect 1324 -168 1326 -156
rect 1339 -161 1341 -145
rect 1368 -157 1370 -144
rect 1455 -152 1457 -127
rect 1471 -140 1473 -137
rect 1486 -140 1488 -137
rect 1515 -140 1517 -137
rect 1471 -152 1473 -145
rect 1455 -156 1473 -152
rect 1363 -159 1370 -157
rect 1329 -164 1330 -161
rect 1334 -164 1341 -161
rect 1368 -164 1370 -159
rect 1339 -168 1341 -164
rect 1471 -168 1473 -156
rect 1486 -161 1488 -145
rect 1515 -157 1517 -144
rect 1594 -152 1596 -127
rect 1610 -140 1612 -137
rect 1625 -140 1627 -137
rect 1654 -140 1656 -137
rect 1610 -152 1612 -145
rect 1594 -156 1612 -152
rect 1510 -159 1517 -157
rect 1476 -164 1477 -161
rect 1481 -164 1488 -161
rect 1515 -164 1517 -159
rect 1486 -168 1488 -164
rect 1610 -168 1612 -156
rect 1625 -161 1627 -145
rect 1654 -157 1656 -144
rect 1718 -152 1720 -127
rect 1734 -140 1736 -137
rect 1749 -140 1751 -137
rect 1778 -140 1780 -137
rect 1734 -152 1736 -145
rect 1718 -156 1736 -152
rect 1649 -159 1656 -157
rect 1615 -164 1616 -161
rect 1620 -164 1627 -161
rect 1654 -164 1656 -159
rect 1625 -168 1627 -164
rect 1734 -168 1736 -156
rect 1749 -161 1751 -145
rect 1778 -157 1780 -144
rect 1773 -159 1780 -157
rect 1739 -164 1740 -161
rect 1744 -164 1751 -161
rect 1778 -164 1780 -159
rect 1749 -168 1751 -164
rect 585 -171 587 -168
rect 110 -181 112 -178
rect 735 -171 737 -168
rect 873 -171 875 -168
rect 1019 -171 1021 -168
rect 1143 -171 1145 -168
rect 1368 -171 1370 -168
rect 1515 -171 1517 -168
rect 1654 -171 1656 -168
rect 1778 -171 1780 -168
rect 691 -178 693 -175
rect 706 -178 708 -175
rect 829 -178 831 -175
rect 844 -178 846 -175
rect 975 -178 977 -175
rect 990 -178 992 -175
rect 1099 -178 1101 -175
rect 1114 -178 1116 -175
rect 1324 -178 1326 -175
rect 1339 -178 1341 -175
rect 1471 -178 1473 -175
rect 1486 -178 1488 -175
rect 1610 -178 1612 -175
rect 1625 -178 1627 -175
rect 1734 -178 1736 -175
rect 1749 -178 1751 -175
rect 378 -187 380 -184
rect 404 -187 406 -184
rect 431 -187 433 -184
rect 545 -185 547 -182
rect 554 -185 556 -182
rect 378 -201 380 -192
rect 404 -201 406 -192
rect 378 -215 380 -205
rect 404 -215 406 -205
rect 431 -204 433 -191
rect 426 -206 433 -204
rect 431 -211 433 -206
rect 431 -218 433 -215
rect 378 -225 380 -222
rect 404 -225 406 -222
rect 378 -253 380 -250
rect 404 -253 406 -250
rect 431 -253 433 -250
rect 2748 -257 2750 575
rect 3219 540 3221 543
rect 3234 540 3236 543
rect 3249 540 3251 543
rect 3264 540 3266 543
rect 3278 540 3280 543
rect 3304 540 3306 543
rect 3219 505 3221 530
rect 3234 505 3236 530
rect 3249 505 3251 530
rect 3264 505 3266 530
rect 3278 505 3280 530
rect 3304 514 3306 530
rect 3321 510 3561 514
rect 3304 505 3306 510
rect 2973 480 2975 483
rect 2973 463 2975 476
rect 3219 464 3221 495
rect 3234 476 3236 495
rect 3249 476 3251 495
rect 3264 476 3266 495
rect 3278 476 3280 495
rect 3304 492 3306 495
rect 378 -267 380 -258
rect 404 -267 406 -258
rect 378 -281 380 -271
rect 404 -281 406 -271
rect 431 -270 433 -257
rect 570 -259 2750 -257
rect 2837 461 2975 463
rect 570 -269 574 -259
rect 426 -272 433 -270
rect 431 -277 433 -272
rect 442 -273 574 -269
rect 686 -273 688 -270
rect 701 -273 703 -270
rect 730 -273 732 -270
rect 431 -284 433 -281
rect 570 -285 574 -273
rect 686 -285 688 -278
rect 378 -291 380 -288
rect 404 -291 406 -288
rect 570 -289 688 -285
rect 686 -301 688 -289
rect 701 -294 703 -278
rect 730 -290 732 -277
rect 807 -285 809 -259
rect 824 -273 826 -270
rect 839 -273 841 -270
rect 868 -273 870 -270
rect 824 -285 826 -278
rect 807 -289 826 -285
rect 725 -292 732 -290
rect 696 -297 703 -294
rect 730 -297 732 -292
rect 701 -301 703 -297
rect 730 -304 732 -301
rect 686 -311 688 -308
rect 701 -311 703 -308
rect 378 -319 380 -316
rect 404 -319 406 -316
rect 431 -319 433 -316
rect 378 -333 380 -324
rect 404 -333 406 -324
rect 378 -347 380 -337
rect 404 -347 406 -337
rect 431 -336 433 -323
rect 426 -338 433 -336
rect 431 -343 433 -338
rect 443 -339 467 -335
rect 431 -350 433 -347
rect 378 -357 380 -354
rect 404 -357 406 -354
rect 463 -390 467 -339
rect 747 -383 749 -293
rect 824 -301 826 -289
rect 839 -294 841 -278
rect 868 -290 870 -277
rect 952 -285 954 -259
rect 970 -273 972 -270
rect 985 -273 987 -270
rect 1014 -273 1016 -270
rect 970 -285 972 -278
rect 952 -289 972 -285
rect 863 -292 870 -290
rect 829 -297 830 -294
rect 834 -297 841 -294
rect 868 -297 870 -292
rect 839 -301 841 -297
rect 868 -304 870 -301
rect 824 -311 826 -308
rect 839 -311 841 -308
rect 885 -378 887 -293
rect 970 -301 972 -289
rect 985 -294 987 -278
rect 1014 -290 1016 -277
rect 1076 -285 1078 -259
rect 1094 -273 1096 -270
rect 1109 -273 1111 -270
rect 1138 -273 1140 -270
rect 1094 -285 1096 -278
rect 1076 -289 1096 -285
rect 1009 -292 1016 -290
rect 975 -297 976 -294
rect 980 -297 987 -294
rect 1014 -297 1016 -292
rect 985 -301 987 -297
rect 1014 -304 1016 -301
rect 970 -311 972 -308
rect 985 -311 987 -308
rect 1028 -373 1030 -293
rect 1094 -301 1096 -289
rect 1109 -294 1111 -278
rect 1138 -290 1140 -277
rect 1303 -285 1305 -259
rect 1319 -273 1321 -270
rect 1334 -273 1336 -270
rect 1363 -273 1365 -270
rect 1319 -285 1321 -278
rect 1303 -289 1321 -285
rect 1133 -292 1140 -290
rect 1099 -297 1100 -294
rect 1104 -297 1111 -294
rect 1138 -297 1140 -292
rect 1109 -301 1111 -297
rect 1138 -304 1140 -301
rect 1094 -311 1096 -308
rect 1109 -311 1111 -308
rect 1152 -368 1154 -293
rect 1319 -301 1321 -289
rect 1334 -294 1336 -278
rect 1363 -290 1365 -277
rect 1449 -285 1451 -259
rect 1466 -273 1468 -270
rect 1481 -273 1483 -270
rect 1510 -273 1512 -270
rect 1466 -285 1468 -278
rect 1449 -289 1468 -285
rect 1358 -292 1365 -290
rect 1324 -297 1325 -294
rect 1329 -297 1336 -294
rect 1363 -297 1365 -292
rect 1334 -301 1336 -297
rect 1363 -304 1365 -301
rect 1319 -311 1321 -308
rect 1334 -311 1336 -308
rect 1379 -363 1381 -293
rect 1466 -301 1468 -289
rect 1481 -294 1483 -278
rect 1510 -290 1512 -277
rect 1588 -285 1590 -259
rect 1605 -273 1607 -270
rect 1620 -273 1622 -270
rect 1649 -273 1651 -270
rect 1605 -285 1607 -278
rect 1588 -289 1607 -285
rect 1505 -292 1512 -290
rect 1471 -297 1472 -294
rect 1476 -297 1483 -294
rect 1510 -297 1512 -292
rect 1481 -301 1483 -297
rect 1510 -304 1512 -301
rect 1466 -311 1468 -308
rect 1481 -311 1483 -308
rect 1528 -358 1530 -293
rect 1605 -301 1607 -289
rect 1620 -294 1622 -278
rect 1649 -290 1651 -277
rect 1711 -285 1713 -259
rect 1729 -273 1731 -270
rect 1744 -273 1746 -270
rect 1773 -273 1775 -270
rect 1729 -285 1731 -278
rect 1711 -289 1731 -285
rect 1644 -292 1651 -290
rect 1610 -297 1611 -294
rect 1615 -297 1622 -294
rect 1649 -297 1651 -292
rect 1620 -301 1622 -297
rect 1649 -304 1651 -301
rect 1605 -311 1607 -308
rect 1620 -311 1622 -308
rect 1665 -353 1667 -295
rect 1729 -301 1731 -289
rect 1744 -294 1746 -278
rect 1773 -290 1775 -277
rect 1768 -292 1775 -290
rect 1734 -297 1735 -294
rect 1739 -297 1746 -294
rect 1773 -297 1775 -292
rect 1744 -301 1746 -297
rect 1773 -304 1775 -301
rect 1729 -311 1731 -308
rect 1744 -311 1746 -308
rect 2726 -349 2735 -347
rect 2726 -353 2728 -349
rect 1665 -355 2728 -353
rect 1528 -360 2810 -358
rect 1379 -365 2793 -363
rect 1152 -370 2772 -368
rect 1028 -375 2763 -373
rect 885 -380 2755 -378
rect 747 -385 2726 -383
rect 463 -392 1710 -390
rect 664 -424 667 -392
rect 682 -412 684 -409
rect 697 -412 699 -409
rect 726 -412 728 -409
rect 682 -424 684 -417
rect 664 -428 684 -424
rect 682 -440 684 -428
rect 697 -433 699 -417
rect 726 -429 728 -416
rect 803 -424 805 -392
rect 820 -412 822 -409
rect 835 -412 837 -409
rect 864 -412 866 -409
rect 820 -424 822 -417
rect 803 -428 822 -424
rect 721 -431 728 -429
rect 687 -436 688 -433
rect 692 -436 699 -433
rect 726 -436 728 -431
rect 738 -432 743 -428
rect 697 -440 699 -436
rect 726 -443 728 -440
rect 682 -450 684 -447
rect 697 -450 699 -447
rect 741 -814 743 -432
rect 820 -440 822 -428
rect 835 -433 837 -417
rect 864 -429 866 -416
rect 949 -424 951 -392
rect 966 -412 968 -409
rect 981 -412 983 -409
rect 1010 -412 1012 -409
rect 966 -424 968 -417
rect 949 -428 968 -424
rect 859 -431 866 -429
rect 825 -436 826 -433
rect 830 -436 837 -433
rect 864 -436 866 -431
rect 835 -440 837 -436
rect 966 -440 968 -428
rect 981 -433 983 -417
rect 1010 -429 1012 -416
rect 1073 -424 1075 -392
rect 1090 -412 1092 -409
rect 1105 -412 1107 -409
rect 1134 -412 1136 -409
rect 1090 -424 1092 -417
rect 1073 -428 1092 -424
rect 1005 -431 1012 -429
rect 971 -436 972 -433
rect 976 -436 983 -433
rect 1010 -436 1012 -431
rect 981 -440 983 -436
rect 1090 -440 1092 -428
rect 1105 -433 1107 -417
rect 1134 -429 1136 -416
rect 1299 -424 1301 -392
rect 1315 -412 1317 -409
rect 1330 -412 1332 -409
rect 1359 -412 1361 -409
rect 1315 -424 1317 -417
rect 1299 -428 1317 -424
rect 1129 -431 1136 -429
rect 1095 -436 1096 -433
rect 1100 -436 1107 -433
rect 1134 -436 1136 -431
rect 1105 -440 1107 -436
rect 1315 -440 1317 -428
rect 1330 -433 1332 -417
rect 1359 -429 1361 -416
rect 1444 -424 1446 -392
rect 1462 -412 1464 -409
rect 1477 -412 1479 -409
rect 1506 -412 1508 -409
rect 1462 -424 1464 -417
rect 1444 -428 1464 -424
rect 1354 -431 1361 -429
rect 1325 -436 1332 -433
rect 1359 -436 1361 -431
rect 1330 -440 1332 -436
rect 864 -443 866 -440
rect 1010 -443 1012 -440
rect 1134 -443 1136 -440
rect 1359 -443 1361 -440
rect 820 -450 822 -447
rect 835 -450 837 -447
rect 966 -450 968 -447
rect 981 -450 983 -447
rect 1090 -450 1092 -447
rect 1105 -450 1107 -447
rect 1315 -450 1317 -447
rect 1330 -450 1332 -447
rect 1371 -790 1373 -428
rect 1462 -440 1464 -428
rect 1477 -433 1479 -417
rect 1506 -429 1508 -416
rect 1584 -424 1586 -392
rect 1601 -412 1603 -409
rect 1616 -412 1618 -409
rect 1645 -412 1647 -409
rect 1601 -424 1603 -417
rect 1584 -428 1603 -424
rect 1501 -431 1508 -429
rect 1467 -436 1468 -433
rect 1472 -436 1479 -433
rect 1506 -436 1508 -431
rect 1518 -432 1521 -428
rect 1477 -440 1479 -436
rect 1506 -443 1508 -440
rect 1462 -450 1464 -447
rect 1477 -450 1479 -447
rect 1519 -680 1521 -432
rect 1601 -440 1603 -428
rect 1616 -433 1618 -417
rect 1645 -429 1647 -416
rect 1708 -424 1710 -392
rect 1725 -412 1727 -409
rect 1740 -412 1742 -409
rect 1769 -412 1771 -409
rect 1725 -424 1727 -417
rect 1708 -428 1727 -424
rect 1640 -431 1647 -429
rect 1606 -436 1607 -433
rect 1611 -436 1618 -433
rect 1645 -436 1647 -431
rect 1657 -432 1660 -428
rect 1616 -440 1618 -436
rect 1645 -443 1647 -440
rect 1601 -450 1603 -447
rect 1616 -450 1618 -447
rect 1658 -559 1660 -432
rect 1725 -440 1727 -428
rect 1740 -433 1742 -417
rect 1769 -429 1771 -416
rect 1764 -431 1771 -429
rect 1730 -436 1731 -433
rect 1735 -436 1742 -433
rect 1769 -436 1771 -431
rect 1740 -440 1742 -436
rect 1769 -443 1771 -440
rect 1725 -450 1727 -447
rect 1740 -450 1742 -447
rect 1781 -468 1783 -428
rect 2724 -438 2726 -385
rect 1841 -456 1843 -453
rect 1856 -456 1858 -453
rect 1885 -456 1887 -453
rect 1841 -468 1843 -461
rect 1781 -472 1843 -468
rect 1841 -484 1843 -472
rect 1856 -477 1858 -461
rect 1885 -473 1887 -460
rect 1880 -475 1887 -473
rect 1846 -480 1847 -477
rect 1851 -480 1858 -477
rect 1885 -480 1887 -475
rect 1856 -484 1858 -480
rect 1885 -487 1887 -484
rect 1841 -494 1843 -491
rect 1856 -494 1858 -491
rect 2753 -529 2755 -380
rect 2761 -386 2763 -375
rect 2769 -375 2772 -370
rect 2761 -388 2784 -386
rect 1658 -561 1826 -559
rect 1841 -561 1843 -558
rect 1856 -561 1858 -558
rect 1885 -561 1887 -558
rect 1824 -573 1826 -561
rect 2782 -563 2784 -388
rect 2791 -393 2793 -365
rect 2807 -385 2810 -360
rect 2837 -371 2839 461
rect 2973 456 2975 461
rect 2985 460 3221 464
rect 2973 449 2975 452
rect 3350 440 3352 443
rect 3365 440 3367 443
rect 3385 440 3387 443
rect 3395 440 3397 443
rect 3421 440 3423 443
rect 3558 432 3561 510
rect 3668 487 3670 490
rect 3680 487 3682 490
rect 3695 487 3697 490
rect 3705 487 3707 490
rect 3728 487 3730 490
rect 3668 457 3670 480
rect 3680 457 3682 480
rect 3695 457 3697 480
rect 3705 457 3707 480
rect 3728 465 3730 480
rect 3728 457 3730 461
rect 3668 432 3670 450
rect 2975 414 2977 417
rect 2975 397 2977 410
rect 3350 405 3352 430
rect 3365 405 3367 430
rect 3385 405 3387 430
rect 3395 405 3397 430
rect 3421 414 3423 430
rect 3558 429 3670 432
rect 3680 414 3682 450
rect 3438 410 3682 414
rect 3421 405 3423 410
rect 2844 395 2977 397
rect 2844 -223 2846 395
rect 2975 390 2977 395
rect 2995 394 3320 398
rect 3488 402 3490 405
rect 3503 402 3505 405
rect 3523 402 3525 405
rect 3547 402 3549 405
rect 2975 383 2977 386
rect 3318 376 3320 394
rect 3350 376 3352 395
rect 3318 374 3352 376
rect 2978 347 2980 350
rect 2978 330 2980 343
rect 2851 328 2980 330
rect 2851 -69 2853 328
rect 2978 323 2980 328
rect 2978 316 2980 319
rect 2978 280 2980 283
rect 2978 263 2980 276
rect 2868 261 2980 263
rect 2868 92 2870 261
rect 2978 256 2980 261
rect 2978 249 2980 252
rect 2996 175 2998 178
rect 2881 168 2917 170
rect 2868 89 2873 92
rect 2881 83 2883 168
rect 2896 139 2898 142
rect 2915 139 2917 168
rect 2996 158 2998 171
rect 2991 156 2998 158
rect 2996 151 2998 156
rect 2996 144 2998 147
rect 2940 139 2942 142
rect 2959 139 2961 142
rect 2896 122 2898 134
rect 2915 131 2917 134
rect 2940 122 2942 134
rect 2896 120 2917 122
rect 2896 108 2898 111
rect 2915 108 2917 120
rect 2941 118 2942 122
rect 2940 108 2942 118
rect 2959 108 2961 134
rect 2970 119 2976 121
rect 2896 83 2898 103
rect 2915 92 2917 103
rect 2940 100 2942 103
rect 2959 92 2961 103
rect 2919 90 2961 92
rect 2974 83 2976 119
rect 2881 81 2976 83
rect 2998 14 3000 17
rect 2883 7 2919 9
rect 2851 -72 2875 -69
rect 2883 -78 2885 7
rect 2898 -22 2900 -19
rect 2917 -22 2919 7
rect 2998 -3 3000 10
rect 2993 -5 3000 -3
rect 2998 -10 3000 -5
rect 2998 -17 3000 -14
rect 2942 -22 2944 -19
rect 2961 -22 2963 -19
rect 2898 -39 2900 -27
rect 2917 -30 2919 -27
rect 2942 -39 2944 -27
rect 2898 -41 2919 -39
rect 2898 -53 2900 -50
rect 2917 -53 2919 -41
rect 2943 -43 2944 -39
rect 2942 -53 2944 -43
rect 2961 -53 2963 -27
rect 2972 -42 2978 -40
rect 2898 -78 2900 -58
rect 2917 -69 2919 -58
rect 2942 -61 2944 -58
rect 2961 -69 2963 -58
rect 2921 -71 2963 -69
rect 2976 -78 2978 -42
rect 2883 -80 2978 -78
rect 3365 -117 3367 395
rect 3385 376 3387 395
rect 3395 375 3397 395
rect 3421 392 3423 395
rect 3488 367 3490 392
rect 3503 367 3505 392
rect 3523 367 3525 392
rect 3547 376 3549 392
rect 3695 376 3697 450
rect 3564 372 3697 376
rect 3547 367 3549 372
rect 3614 357 3616 360
rect 3635 357 3637 360
rect 3661 357 3663 360
rect 3488 338 3490 357
rect 3503 316 3505 357
rect 3523 337 3525 357
rect 3547 354 3549 357
rect 3614 329 3616 352
rect 3635 329 3637 352
rect 3661 340 3663 353
rect 3705 341 3707 450
rect 3728 447 3730 450
rect 3656 338 3663 340
rect 3661 333 3663 338
rect 3672 337 3707 341
rect 3661 326 3663 329
rect 3614 264 3616 322
rect 3635 311 3637 322
rect 3428 260 3616 264
rect 3757 -24 3759 575
rect 3735 -26 3759 -24
rect 3597 -34 3599 -31
rect 3612 -34 3614 -31
rect 3632 -34 3634 -31
rect 3642 -34 3644 -31
rect 3668 -34 3670 -31
rect 3709 -41 3711 -38
rect 3735 -41 3737 -26
rect 3767 -41 3769 -38
rect 3597 -69 3599 -44
rect 3612 -69 3614 -44
rect 3632 -69 3634 -44
rect 3642 -69 3644 -44
rect 3668 -60 3670 -44
rect 3709 -55 3711 -46
rect 3735 -55 3737 -46
rect 3668 -69 3670 -64
rect 3709 -69 3711 -59
rect 3735 -69 3737 -59
rect 3767 -58 3769 -45
rect 3762 -60 3769 -58
rect 3767 -65 3769 -60
rect 3767 -72 3769 -69
rect 3709 -79 3711 -76
rect 3735 -79 3737 -76
rect 3597 -96 3599 -79
rect 3574 -98 3599 -96
rect 3612 -103 3614 -79
rect 3574 -105 3614 -103
rect 3632 -111 3634 -79
rect 3574 -113 3634 -111
rect 2912 -121 3367 -117
rect 3642 -119 3644 -79
rect 3668 -82 3670 -79
rect 3574 -121 3644 -119
rect 2997 -140 2999 -137
rect 2882 -147 2918 -145
rect 2844 -226 2874 -223
rect 2882 -232 2884 -147
rect 2897 -176 2899 -173
rect 2916 -176 2918 -147
rect 2997 -157 2999 -144
rect 2992 -159 2999 -157
rect 2997 -164 2999 -159
rect 2997 -171 2999 -168
rect 2941 -176 2943 -173
rect 2960 -176 2962 -173
rect 2897 -193 2899 -181
rect 2916 -184 2918 -181
rect 2941 -193 2943 -181
rect 2897 -195 2918 -193
rect 2897 -207 2899 -204
rect 2916 -207 2918 -195
rect 2942 -197 2943 -193
rect 2941 -207 2943 -197
rect 2960 -207 2962 -181
rect 2971 -196 2977 -194
rect 2897 -232 2899 -212
rect 2916 -223 2918 -212
rect 2941 -215 2943 -212
rect 2960 -223 2962 -212
rect 2920 -225 2962 -223
rect 2975 -232 2977 -196
rect 2882 -234 2977 -232
rect 2997 -288 2999 -285
rect 2882 -295 2918 -293
rect 2837 -374 2874 -371
rect 2882 -380 2884 -295
rect 2897 -324 2899 -321
rect 2916 -324 2918 -295
rect 2997 -305 2999 -292
rect 3659 -293 3661 -290
rect 3671 -293 3673 -290
rect 3686 -293 3688 -290
rect 3696 -293 3698 -290
rect 3719 -293 3721 -290
rect 2992 -307 2999 -305
rect 2997 -312 2999 -307
rect 2997 -319 2999 -316
rect 2941 -324 2943 -321
rect 2960 -324 2962 -321
rect 3659 -323 3661 -300
rect 3671 -323 3673 -300
rect 3686 -323 3688 -300
rect 3696 -323 3698 -300
rect 3719 -315 3721 -300
rect 3719 -323 3721 -319
rect 2897 -341 2899 -329
rect 2916 -332 2918 -329
rect 2941 -341 2943 -329
rect 2897 -343 2918 -341
rect 2897 -355 2899 -352
rect 2916 -355 2918 -343
rect 2942 -345 2943 -341
rect 2941 -355 2943 -345
rect 2960 -355 2962 -329
rect 2971 -344 2977 -342
rect 2897 -380 2899 -360
rect 2916 -371 2918 -360
rect 2941 -363 2943 -360
rect 2960 -371 2962 -360
rect 2920 -373 2962 -371
rect 2975 -380 2977 -344
rect 3434 -349 3436 -346
rect 3449 -349 3451 -346
rect 3464 -349 3466 -346
rect 3479 -349 3481 -346
rect 3493 -349 3495 -346
rect 3519 -349 3521 -346
rect 2882 -382 2977 -380
rect 3434 -384 3436 -359
rect 3449 -384 3451 -359
rect 3464 -384 3466 -359
rect 3479 -384 3481 -359
rect 3493 -384 3495 -359
rect 3519 -375 3521 -359
rect 3659 -375 3661 -330
rect 3536 -379 3661 -375
rect 3519 -384 3521 -379
rect 2807 -388 2852 -385
rect 2907 -393 2909 -391
rect 2791 -395 2909 -393
rect 2973 -415 2975 -412
rect 3434 -414 3436 -394
rect 3449 -414 3451 -394
rect 3464 -414 3466 -394
rect 3479 -413 3481 -394
rect 3493 -413 3495 -394
rect 3519 -397 3521 -394
rect 3212 -417 3436 -414
rect 2973 -432 2975 -419
rect 3212 -431 3217 -417
rect 2955 -434 2975 -432
rect 2960 -439 2962 -434
rect 2973 -439 2975 -434
rect 3039 -435 3217 -431
rect 3302 -433 3304 -430
rect 3317 -433 3319 -430
rect 3337 -433 3339 -430
rect 3347 -433 3349 -430
rect 3373 -433 3375 -430
rect 2801 -442 2962 -439
rect 2973 -446 2975 -443
rect 3302 -468 3304 -443
rect 3317 -468 3319 -443
rect 3337 -468 3339 -443
rect 3347 -468 3349 -443
rect 3373 -459 3375 -443
rect 3671 -459 3673 -330
rect 3686 -343 3688 -330
rect 3390 -463 3673 -459
rect 3373 -468 3375 -463
rect 2975 -481 2977 -478
rect 2975 -498 2977 -485
rect 3302 -497 3304 -478
rect 3317 -497 3319 -478
rect 3337 -496 3339 -478
rect 3347 -496 3349 -478
rect 3373 -481 3375 -478
rect 2955 -500 2977 -498
rect 2975 -505 2977 -500
rect 2996 -500 3304 -497
rect 3161 -508 3163 -505
rect 3176 -508 3178 -505
rect 3196 -508 3198 -505
rect 3220 -508 3222 -505
rect 2975 -512 2977 -509
rect 3161 -543 3163 -518
rect 3176 -543 3178 -518
rect 3196 -543 3198 -518
rect 3220 -534 3222 -518
rect 3220 -543 3222 -538
rect 2978 -548 2980 -545
rect 1841 -573 1843 -566
rect 1824 -577 1843 -573
rect 1841 -589 1843 -577
rect 1856 -582 1858 -566
rect 1885 -578 1887 -565
rect 2782 -566 2846 -563
rect 2978 -565 2980 -552
rect 2955 -567 2980 -565
rect 2978 -572 2980 -567
rect 2990 -568 3143 -564
rect 3140 -574 3143 -568
rect 3161 -574 3163 -553
rect 3176 -572 3178 -553
rect 1880 -580 1887 -578
rect 2978 -579 2980 -576
rect 3140 -577 3163 -574
rect 3196 -573 3198 -553
rect 3220 -556 3222 -553
rect 1846 -585 1847 -582
rect 1851 -585 1858 -582
rect 1885 -585 1887 -580
rect 1856 -589 1858 -585
rect 3063 -587 3065 -584
rect 3084 -587 3086 -584
rect 3110 -587 3112 -584
rect 1885 -592 1887 -589
rect 1841 -599 1843 -596
rect 1856 -599 1858 -596
rect 2978 -615 2980 -612
rect 3063 -615 3065 -592
rect 3084 -615 3086 -592
rect 3110 -604 3112 -591
rect 3696 -603 3698 -330
rect 3719 -333 3721 -330
rect 3105 -606 3112 -604
rect 3110 -611 3112 -606
rect 3121 -607 3698 -603
rect 2978 -632 2980 -619
rect 3110 -618 3112 -615
rect 3063 -631 3065 -622
rect 2955 -634 2980 -632
rect 2978 -639 2980 -634
rect 2991 -635 3065 -631
rect 3084 -635 3086 -622
rect 2978 -646 2980 -643
rect 1519 -682 1823 -680
rect 1821 -695 1823 -682
rect 1841 -683 1843 -680
rect 1856 -683 1858 -680
rect 1885 -683 1887 -680
rect 1841 -695 1843 -688
rect 1821 -699 1843 -695
rect 1841 -711 1843 -699
rect 1856 -704 1858 -688
rect 1885 -700 1887 -687
rect 1880 -702 1887 -700
rect 1846 -707 1847 -704
rect 1851 -707 1858 -704
rect 1885 -707 1887 -702
rect 1856 -711 1858 -707
rect 1885 -714 1887 -711
rect 1841 -721 1843 -718
rect 1856 -721 1858 -718
rect 1841 -790 1843 -787
rect 1856 -790 1858 -787
rect 1885 -790 1887 -787
rect 1371 -792 1825 -790
rect 1823 -802 1825 -792
rect 1841 -802 1843 -795
rect 1823 -806 1843 -802
rect 1811 -814 1833 -811
rect 741 -815 1833 -814
rect 741 -816 1813 -815
rect 1841 -818 1843 -806
rect 1856 -811 1858 -795
rect 1885 -807 1887 -794
rect 1880 -809 1887 -807
rect 1846 -814 1847 -811
rect 1851 -814 1858 -811
rect 1885 -814 1887 -809
rect 1856 -818 1858 -814
rect 1885 -821 1887 -818
rect 1841 -828 1843 -825
rect 1856 -828 1858 -825
<< polycontact >>
rect 2139 915 2143 919
rect 2168 915 2172 919
rect 2117 885 2121 889
rect 2276 911 2280 915
rect 2305 911 2309 915
rect 2252 882 2256 886
rect 2127 848 2131 852
rect 2164 844 2168 848
rect 2340 854 2344 858
rect 2135 839 2139 843
rect 2212 838 2216 842
rect 2229 838 2233 842
rect 2266 834 2270 838
rect 2384 853 2388 857
rect 2359 847 2363 851
rect 2401 853 2405 857
rect 2237 829 2241 833
rect 2212 802 2216 806
rect 2137 639 2141 643
rect 2166 639 2170 643
rect 2115 609 2119 613
rect 2274 635 2278 639
rect 2303 635 2307 639
rect 2250 606 2254 610
rect 2125 572 2129 576
rect 2162 568 2166 572
rect 2338 578 2342 582
rect 2133 563 2137 567
rect 2210 562 2214 566
rect 2227 562 2231 566
rect 2264 558 2268 562
rect 2382 577 2386 581
rect 2357 571 2361 575
rect 2235 553 2239 557
rect 2134 360 2138 364
rect 2163 360 2167 364
rect 2112 330 2116 334
rect 2271 356 2275 360
rect 2300 356 2304 360
rect 2247 327 2251 331
rect 2122 293 2126 297
rect 2159 289 2163 293
rect 2335 299 2339 303
rect 2130 284 2134 288
rect 2207 283 2211 287
rect 2224 283 2228 287
rect 2261 279 2265 283
rect 2379 298 2383 302
rect 2354 292 2358 296
rect 2396 298 2400 302
rect 2232 274 2236 278
rect 2207 247 2211 251
rect 1474 14 1478 18
rect 1503 14 1507 18
rect 1452 -16 1456 -12
rect 1623 12 1627 16
rect 1652 12 1656 16
rect 1601 -18 1605 -14
rect 1775 11 1779 15
rect 1804 11 1808 15
rect 1753 -19 1757 -15
rect 2137 75 2141 79
rect 2166 75 2170 79
rect 2115 45 2119 49
rect 2274 71 2278 75
rect 2303 71 2307 75
rect 2250 42 2254 46
rect 1926 10 1930 14
rect 1955 10 1959 14
rect 1904 -20 1908 -16
rect 2125 8 2129 12
rect 2162 4 2166 8
rect 2338 14 2342 18
rect 2133 -1 2137 3
rect 2210 -2 2214 2
rect 2227 -2 2231 2
rect 2264 -6 2268 -2
rect 2382 13 2386 17
rect 2357 7 2361 11
rect 2235 -11 2239 -7
rect 101 -115 105 -111
rect 376 -136 380 -132
rect 402 -136 406 -132
rect 422 -138 426 -134
rect 101 -170 105 -166
rect 1198 -81 1202 -77
rect 1241 -76 1245 -72
rect 1212 -81 1216 -77
rect 532 -159 536 -155
rect 517 -167 521 -163
rect 576 -160 580 -156
rect 551 -166 555 -162
rect 593 -160 597 -156
rect 726 -160 730 -156
rect 697 -165 701 -161
rect 864 -160 868 -156
rect 835 -165 839 -161
rect 1010 -160 1014 -156
rect 981 -165 985 -161
rect 1134 -160 1138 -156
rect 1105 -165 1109 -161
rect 1359 -160 1363 -156
rect 1330 -165 1334 -161
rect 1506 -160 1510 -156
rect 1477 -165 1481 -161
rect 1645 -160 1649 -156
rect 1616 -165 1620 -161
rect 1769 -160 1773 -156
rect 1740 -165 1744 -161
rect 376 -205 380 -201
rect 402 -205 406 -201
rect 422 -207 426 -203
rect 3302 510 3306 514
rect 3317 510 3321 514
rect 3233 472 3237 476
rect 3248 472 3252 476
rect 3263 472 3267 476
rect 3277 472 3281 476
rect 376 -271 380 -267
rect 402 -271 406 -267
rect 422 -273 426 -269
rect 438 -273 442 -269
rect 721 -293 725 -289
rect 692 -298 696 -294
rect 745 -293 749 -289
rect 376 -337 380 -333
rect 402 -337 406 -333
rect 422 -339 426 -335
rect 439 -339 443 -335
rect 859 -293 863 -289
rect 830 -298 834 -294
rect 884 -293 888 -289
rect 1005 -293 1009 -289
rect 976 -298 980 -294
rect 1027 -293 1031 -289
rect 1129 -293 1133 -289
rect 1100 -298 1104 -294
rect 1151 -293 1155 -289
rect 1354 -293 1358 -289
rect 1325 -298 1329 -294
rect 1378 -293 1382 -289
rect 1501 -293 1505 -289
rect 1472 -298 1476 -294
rect 1527 -293 1531 -289
rect 1640 -293 1644 -289
rect 1611 -298 1615 -294
rect 1664 -295 1668 -291
rect 1764 -293 1768 -289
rect 1735 -298 1739 -294
rect 2735 -350 2739 -346
rect 717 -432 721 -428
rect 688 -437 692 -433
rect 734 -432 738 -428
rect 855 -432 859 -428
rect 826 -437 830 -433
rect 1001 -432 1005 -428
rect 972 -437 976 -433
rect 1125 -432 1129 -428
rect 1096 -437 1100 -433
rect 1350 -432 1354 -428
rect 1321 -437 1325 -433
rect 1367 -432 1371 -428
rect 1497 -432 1501 -428
rect 1468 -437 1472 -433
rect 1514 -432 1518 -428
rect 1636 -432 1640 -428
rect 1607 -437 1611 -433
rect 1653 -432 1657 -428
rect 1760 -432 1764 -428
rect 1731 -437 1735 -433
rect 1777 -432 1781 -428
rect 2724 -442 2728 -438
rect 1876 -476 1880 -472
rect 1847 -481 1851 -477
rect 2769 -379 2773 -375
rect 2752 -533 2756 -529
rect 2981 460 2985 464
rect 3726 461 3730 465
rect 3419 410 3423 414
rect 3434 410 3438 414
rect 2991 394 2995 398
rect 2873 88 2877 92
rect 2987 155 2991 159
rect 2937 118 2941 122
rect 2966 118 2970 122
rect 2915 88 2919 92
rect 2875 -73 2879 -69
rect 2989 -6 2993 -2
rect 2939 -43 2943 -39
rect 2968 -43 2972 -39
rect 2917 -73 2921 -69
rect 3384 372 3388 376
rect 3394 371 3398 375
rect 3545 372 3549 376
rect 3560 372 3564 376
rect 3487 334 3491 338
rect 3522 333 3526 337
rect 3652 337 3656 341
rect 3668 337 3672 341
rect 3502 312 3506 316
rect 3634 307 3638 311
rect 3424 260 3428 264
rect 3707 -59 3711 -55
rect 3733 -59 3737 -55
rect 3666 -64 3670 -60
rect 3758 -61 3762 -57
rect 3570 -98 3574 -94
rect 3570 -106 3574 -102
rect 3570 -114 3574 -110
rect 2908 -121 2912 -117
rect 3570 -122 3574 -118
rect 2874 -227 2878 -223
rect 2988 -160 2992 -156
rect 2938 -197 2942 -193
rect 2967 -197 2971 -193
rect 2916 -227 2920 -223
rect 2874 -375 2878 -371
rect 2988 -308 2992 -304
rect 3717 -319 3721 -315
rect 2938 -345 2942 -341
rect 2967 -345 2971 -341
rect 2916 -375 2920 -371
rect 3517 -379 3521 -375
rect 3532 -379 3536 -375
rect 2852 -389 2856 -385
rect 2907 -391 2911 -387
rect 2951 -435 2955 -431
rect 3448 -418 3452 -414
rect 3463 -418 3467 -414
rect 3478 -417 3482 -413
rect 3492 -417 3496 -413
rect 3035 -435 3039 -431
rect 2797 -443 2801 -439
rect 3685 -347 3689 -343
rect 3371 -463 3375 -459
rect 3386 -463 3390 -459
rect 2951 -501 2955 -497
rect 2992 -501 2996 -497
rect 3316 -501 3320 -497
rect 3336 -500 3340 -496
rect 3346 -500 3350 -496
rect 3218 -538 3222 -534
rect 1876 -581 1880 -577
rect 2846 -566 2850 -562
rect 2951 -568 2955 -564
rect 2986 -568 2990 -564
rect 3175 -576 3179 -572
rect 3195 -577 3199 -573
rect 1847 -586 1851 -582
rect 3101 -607 3105 -603
rect 3117 -607 3121 -603
rect 2951 -635 2955 -631
rect 2987 -635 2991 -631
rect 3083 -639 3087 -635
rect 1876 -703 1880 -699
rect 1847 -708 1851 -704
rect 1833 -815 1837 -811
rect 1876 -810 1880 -806
rect 1847 -815 1851 -811
<< metal1 >>
rect 51 1053 2471 1083
rect 53 994 69 1053
rect 53 -70 70 994
rect 2182 967 2278 970
rect 2093 959 2133 963
rect 2093 935 2097 959
rect 2093 918 2097 931
rect 2071 915 2097 918
rect 2071 882 2074 915
rect 2093 904 2097 915
rect 2102 952 2120 956
rect 2102 935 2106 952
rect 2121 935 2125 951
rect 2102 904 2106 931
rect 2112 904 2116 931
rect 2121 904 2125 931
rect 2129 919 2133 959
rect 2182 951 2185 967
rect 2137 947 2185 951
rect 2137 935 2141 947
rect 2156 935 2160 947
rect 2129 915 2139 919
rect 2146 911 2150 931
rect 2129 907 2150 911
rect 2112 897 2116 900
rect 2129 897 2133 907
rect 2146 904 2150 907
rect 2165 919 2169 931
rect 2165 915 2168 919
rect 2165 904 2169 915
rect 2112 893 2133 897
rect 2137 897 2141 900
rect 2156 897 2160 900
rect 2137 893 2155 897
rect 2072 876 2074 882
rect 2071 843 2074 876
rect 2077 886 2117 889
rect 2077 867 2080 886
rect 2182 873 2185 947
rect 2230 955 2270 959
rect 2230 931 2234 955
rect 2230 914 2234 927
rect 2216 911 2234 914
rect 2230 900 2234 911
rect 2239 948 2262 952
rect 2239 931 2243 948
rect 2258 931 2262 948
rect 2239 900 2243 927
rect 2249 900 2253 927
rect 2258 900 2262 927
rect 2266 915 2270 955
rect 2274 947 2278 967
rect 2325 947 2332 1053
rect 2274 943 2337 947
rect 2274 931 2278 943
rect 2293 931 2297 943
rect 2266 911 2276 915
rect 2283 907 2287 927
rect 2266 903 2287 907
rect 2249 893 2253 896
rect 2266 893 2270 903
rect 2283 900 2287 903
rect 2302 915 2306 927
rect 2302 911 2305 915
rect 2302 900 2306 911
rect 2249 889 2270 893
rect 2274 893 2278 896
rect 2293 893 2297 896
rect 2274 889 2297 893
rect 2216 882 2252 885
rect 2274 879 2277 889
rect 2193 876 2277 879
rect 2117 869 2202 873
rect 2123 863 2127 869
rect 2077 852 2080 862
rect 2077 848 2127 852
rect 2135 850 2139 860
rect 2149 863 2153 869
rect 2168 864 2171 869
rect 2199 863 2202 869
rect 2135 848 2162 850
rect 2176 848 2179 860
rect 2199 859 2289 863
rect 2225 853 2229 859
rect 2135 847 2164 848
rect 2159 844 2164 847
rect 2176 844 2195 848
rect 2159 843 2162 844
rect 2071 839 2135 843
rect 2149 839 2162 843
rect 2176 840 2179 844
rect 2123 822 2127 832
rect 2149 833 2153 839
rect 2169 825 2172 836
rect 2123 820 2169 822
rect 2123 819 2172 820
rect 2192 814 2195 844
rect 2212 842 2216 850
rect 2216 838 2229 842
rect 2237 840 2241 850
rect 2251 853 2255 859
rect 2270 854 2273 859
rect 2237 838 2264 840
rect 2278 838 2281 850
rect 2237 837 2266 838
rect 2261 834 2266 837
rect 2278 834 2284 838
rect 2261 833 2264 834
rect 2227 829 2237 833
rect 2251 829 2264 833
rect 2278 830 2281 834
rect 2225 812 2229 822
rect 2251 823 2255 829
rect 2271 812 2274 826
rect 2294 825 2297 889
rect 2334 882 2337 943
rect 2334 879 2407 882
rect 2345 873 2349 879
rect 2388 873 2391 879
rect 2338 854 2340 858
rect 2368 855 2372 864
rect 2396 857 2399 869
rect 2379 855 2384 857
rect 2366 853 2384 855
rect 2396 853 2401 857
rect 2366 851 2382 853
rect 2339 847 2359 850
rect 2366 844 2369 851
rect 2396 849 2399 853
rect 2357 841 2369 844
rect 2357 840 2361 841
rect 2389 840 2392 845
rect 2385 837 2392 840
rect 2345 825 2349 831
rect 2368 825 2372 831
rect 2385 825 2388 837
rect 2294 822 2371 825
rect 2294 812 2297 822
rect 2376 822 2388 825
rect 2225 809 2297 812
rect 2212 794 2216 802
rect 2023 791 2216 794
rect 1260 76 1931 79
rect 1260 -47 1263 76
rect 1477 75 1931 76
rect 1428 58 1468 62
rect 1428 34 1432 58
rect 1428 17 1432 30
rect 1394 14 1432 17
rect 1184 -51 1264 -47
rect 53 -74 136 -70
rect 141 -74 491 -70
rect 91 -86 95 -74
rect 91 -90 124 -86
rect 105 -95 108 -90
rect 366 -97 371 -74
rect 113 -111 116 -99
rect 366 -109 371 -102
rect 487 -109 491 -74
rect 69 -115 101 -111
rect 113 -115 254 -111
rect 86 -131 92 -115
rect 113 -119 116 -115
rect 260 -115 355 -111
rect 366 -112 491 -109
rect 106 -127 109 -123
rect 351 -132 355 -115
rect 372 -119 376 -112
rect 351 -136 376 -132
rect 99 -145 121 -141
rect 105 -150 108 -145
rect 179 -143 341 -139
rect 113 -166 116 -154
rect 179 -166 183 -143
rect 383 -139 387 -122
rect 398 -119 402 -112
rect 420 -113 491 -112
rect 426 -118 429 -113
rect 400 -136 402 -132
rect 409 -139 413 -122
rect 434 -134 437 -122
rect 487 -131 491 -113
rect 1184 -131 1187 -51
rect 1200 -57 1204 -51
rect 1212 -70 1216 -60
rect 1226 -57 1230 -51
rect 1245 -56 1248 -51
rect 1212 -72 1239 -70
rect 1253 -72 1256 -60
rect 1394 -72 1397 14
rect 1428 3 1432 14
rect 1437 51 1456 55
rect 1437 34 1441 51
rect 1456 34 1460 50
rect 1437 3 1441 30
rect 1447 3 1451 30
rect 1456 3 1460 30
rect 1464 18 1468 58
rect 1477 50 1481 75
rect 1577 56 1617 60
rect 1472 46 1495 50
rect 1472 34 1476 46
rect 1491 34 1495 46
rect 1464 14 1474 18
rect 1481 10 1485 30
rect 1464 6 1485 10
rect 1447 -4 1451 -1
rect 1464 -4 1468 6
rect 1481 3 1485 6
rect 1500 18 1504 30
rect 1577 32 1581 56
rect 1500 14 1503 18
rect 1577 15 1581 28
rect 1500 3 1504 14
rect 1447 -8 1468 -4
rect 1535 12 1581 15
rect 1472 -4 1476 -1
rect 1491 -4 1495 -1
rect 1472 -8 1482 -4
rect 1487 -8 1495 -4
rect 1416 -15 1452 -12
rect 1535 -72 1538 12
rect 1577 1 1581 12
rect 1586 52 1609 53
rect 1586 49 1604 52
rect 1586 32 1590 49
rect 1605 32 1609 47
rect 1586 1 1590 28
rect 1596 1 1600 28
rect 1605 1 1609 28
rect 1613 16 1617 56
rect 1626 48 1631 75
rect 1729 55 1769 59
rect 1621 44 1644 48
rect 1621 32 1625 44
rect 1640 32 1644 44
rect 1613 12 1623 16
rect 1630 8 1634 28
rect 1613 4 1634 8
rect 1596 -6 1600 -3
rect 1613 -6 1617 4
rect 1630 1 1634 4
rect 1649 16 1653 28
rect 1729 31 1733 55
rect 1649 12 1652 16
rect 1729 14 1733 27
rect 1649 1 1653 12
rect 1596 -10 1617 -6
rect 1694 11 1733 14
rect 1621 -6 1625 -3
rect 1640 -6 1644 -3
rect 1621 -10 1631 -6
rect 1636 -10 1644 -6
rect 1563 -17 1601 -14
rect 1694 -72 1697 11
rect 1729 0 1733 11
rect 1738 48 1756 52
rect 1738 31 1742 48
rect 1757 31 1761 47
rect 1738 0 1742 27
rect 1748 0 1752 27
rect 1757 0 1761 27
rect 1765 15 1769 55
rect 1777 47 1780 75
rect 1880 54 1920 58
rect 1773 43 1796 47
rect 1773 31 1777 43
rect 1792 31 1796 43
rect 1765 11 1775 15
rect 1782 7 1786 27
rect 1765 3 1786 7
rect 1748 -7 1752 -4
rect 1765 -7 1769 3
rect 1782 0 1786 3
rect 1801 15 1805 27
rect 1880 30 1884 54
rect 1801 11 1804 15
rect 1880 13 1884 26
rect 1801 0 1805 11
rect 1748 -11 1769 -7
rect 1851 10 1884 13
rect 1773 -7 1777 -4
rect 1792 -7 1796 -4
rect 1773 -11 1783 -7
rect 1788 -11 1796 -7
rect 1714 -18 1753 -15
rect 1851 -72 1854 10
rect 1880 -1 1884 10
rect 1889 47 1908 51
rect 1889 30 1893 47
rect 1908 30 1912 46
rect 1889 -1 1893 26
rect 1899 -1 1903 26
rect 1908 -1 1912 26
rect 1916 14 1920 54
rect 1927 46 1931 75
rect 1924 42 1947 46
rect 1924 30 1928 42
rect 1943 30 1947 42
rect 1916 10 1926 14
rect 1933 6 1937 26
rect 1916 2 1937 6
rect 1899 -8 1903 -5
rect 1916 -8 1920 2
rect 1933 -1 1937 2
rect 1952 14 1956 26
rect 1952 10 1955 14
rect 1952 -1 1956 10
rect 1899 -12 1920 -8
rect 1924 -8 1928 -5
rect 1943 -8 1947 -5
rect 1924 -12 1933 -8
rect 1938 -12 1947 -8
rect 1866 -19 1904 -16
rect 2023 -71 2029 791
rect 2180 691 2276 694
rect 2091 683 2131 687
rect 2091 659 2095 683
rect 2091 642 2095 655
rect 2069 639 2095 642
rect 2069 602 2072 639
rect 2091 628 2095 639
rect 2100 676 2118 680
rect 2100 659 2104 676
rect 2119 659 2123 675
rect 2100 628 2104 655
rect 2110 628 2114 655
rect 2119 628 2123 655
rect 2127 643 2131 683
rect 2180 675 2183 691
rect 2135 671 2183 675
rect 2135 659 2139 671
rect 2154 659 2158 671
rect 2127 639 2137 643
rect 2144 635 2148 655
rect 2127 631 2148 635
rect 2110 621 2114 624
rect 2127 621 2131 631
rect 2144 628 2148 631
rect 2163 643 2167 655
rect 2163 639 2166 643
rect 2163 628 2167 639
rect 2110 617 2131 621
rect 2135 621 2139 624
rect 2154 621 2158 624
rect 2135 617 2153 621
rect 2069 567 2072 597
rect 2075 610 2115 613
rect 2075 589 2078 610
rect 2180 597 2183 671
rect 2228 679 2268 683
rect 2228 655 2232 679
rect 2228 638 2232 651
rect 2214 635 2232 638
rect 2228 624 2232 635
rect 2237 672 2260 676
rect 2237 655 2241 672
rect 2256 655 2260 672
rect 2237 624 2241 651
rect 2247 624 2251 651
rect 2256 624 2260 651
rect 2264 639 2268 679
rect 2272 671 2276 691
rect 2272 667 2335 671
rect 2272 655 2276 667
rect 2291 655 2295 667
rect 2264 635 2274 639
rect 2281 631 2285 651
rect 2264 627 2285 631
rect 2247 617 2251 620
rect 2264 617 2268 627
rect 2281 624 2285 627
rect 2300 639 2304 651
rect 2300 635 2303 639
rect 2300 624 2304 635
rect 2247 613 2268 617
rect 2272 617 2276 620
rect 2291 617 2295 620
rect 2272 613 2295 617
rect 2214 606 2250 609
rect 2272 603 2275 613
rect 2191 600 2275 603
rect 2115 593 2200 597
rect 2121 587 2125 593
rect 2075 576 2078 584
rect 2075 572 2125 576
rect 2133 574 2137 584
rect 2147 587 2151 593
rect 2166 588 2169 593
rect 2197 587 2200 593
rect 2133 572 2160 574
rect 2174 572 2177 584
rect 2197 583 2287 587
rect 2223 577 2227 583
rect 2133 571 2162 572
rect 2157 568 2162 571
rect 2174 568 2193 572
rect 2157 567 2160 568
rect 2069 563 2133 567
rect 2147 563 2160 567
rect 2174 564 2177 568
rect 2121 546 2125 556
rect 2147 557 2151 563
rect 2167 549 2170 560
rect 2121 544 2167 546
rect 2121 543 2170 544
rect 2190 538 2193 568
rect 2210 566 2214 574
rect 2214 562 2227 566
rect 2235 564 2239 574
rect 2249 577 2253 583
rect 2268 578 2271 583
rect 2235 562 2262 564
rect 2276 562 2279 574
rect 2235 561 2264 562
rect 2259 558 2264 561
rect 2276 558 2282 562
rect 2259 557 2262 558
rect 2225 553 2235 557
rect 2249 553 2262 557
rect 2276 554 2279 558
rect 2223 536 2227 546
rect 2249 547 2253 553
rect 2269 536 2272 550
rect 2292 549 2295 613
rect 2332 606 2335 667
rect 2463 606 2470 1053
rect 2332 603 2448 606
rect 2343 597 2347 603
rect 2386 597 2389 603
rect 2453 603 2470 606
rect 2336 578 2338 582
rect 2366 579 2370 588
rect 2394 581 2397 593
rect 2377 579 2382 581
rect 2364 577 2382 579
rect 2394 577 2430 581
rect 2364 575 2380 577
rect 2337 571 2357 574
rect 2364 568 2367 575
rect 2394 573 2397 577
rect 2355 565 2367 568
rect 2355 564 2359 565
rect 2387 564 2390 569
rect 2383 561 2390 564
rect 2343 549 2347 555
rect 2366 549 2370 555
rect 2383 549 2386 561
rect 2292 546 2370 549
rect 2292 536 2295 546
rect 2375 546 2386 549
rect 2223 533 2295 536
rect 2177 412 2273 415
rect 2088 404 2128 408
rect 2088 380 2092 404
rect 2088 363 2092 376
rect 2066 360 2092 363
rect 2066 328 2069 360
rect 2088 349 2092 360
rect 2097 397 2115 401
rect 2097 380 2101 397
rect 2116 380 2120 396
rect 2097 349 2101 376
rect 2107 349 2111 376
rect 2116 349 2120 376
rect 2124 364 2128 404
rect 2177 396 2180 412
rect 2132 392 2180 396
rect 2132 380 2136 392
rect 2151 380 2155 392
rect 2124 360 2134 364
rect 2141 356 2145 376
rect 2124 352 2145 356
rect 2107 342 2111 345
rect 2124 342 2128 352
rect 2141 349 2145 352
rect 2160 364 2164 376
rect 2160 360 2163 364
rect 2160 349 2164 360
rect 2107 338 2128 342
rect 2132 342 2136 345
rect 2151 342 2155 345
rect 2132 338 2150 342
rect 2068 323 2069 328
rect 2066 288 2069 323
rect 2072 331 2112 334
rect 2072 313 2075 331
rect 2177 318 2180 392
rect 2225 400 2265 404
rect 2225 376 2229 400
rect 2225 359 2229 372
rect 2211 356 2229 359
rect 2225 345 2229 356
rect 2234 393 2257 397
rect 2234 376 2238 393
rect 2253 376 2257 393
rect 2234 345 2238 372
rect 2244 345 2248 372
rect 2253 345 2257 372
rect 2261 360 2265 400
rect 2269 392 2273 412
rect 2269 388 2332 392
rect 2269 376 2273 388
rect 2288 376 2292 388
rect 2261 356 2271 360
rect 2278 352 2282 372
rect 2261 348 2282 352
rect 2244 338 2248 341
rect 2261 338 2265 348
rect 2278 345 2282 348
rect 2297 360 2301 372
rect 2297 356 2300 360
rect 2297 345 2301 356
rect 2244 334 2265 338
rect 2269 338 2273 341
rect 2288 338 2292 341
rect 2269 334 2292 338
rect 2211 327 2247 330
rect 2269 324 2272 334
rect 2188 321 2272 324
rect 2112 314 2197 318
rect 2118 308 2122 314
rect 2072 297 2075 308
rect 2072 293 2122 297
rect 2130 295 2134 305
rect 2144 308 2148 314
rect 2163 309 2166 314
rect 2194 308 2197 314
rect 2130 293 2157 295
rect 2171 293 2174 305
rect 2194 304 2284 308
rect 2220 298 2224 304
rect 2130 292 2159 293
rect 2154 289 2159 292
rect 2171 289 2190 293
rect 2154 288 2157 289
rect 2066 284 2130 288
rect 2144 284 2157 288
rect 2171 285 2174 289
rect 2118 267 2122 277
rect 2144 278 2148 284
rect 2164 270 2167 281
rect 2118 265 2164 267
rect 2118 264 2167 265
rect 2187 259 2190 289
rect 2207 287 2211 295
rect 2211 283 2224 287
rect 2232 285 2236 295
rect 2246 298 2250 304
rect 2265 299 2268 304
rect 2232 283 2259 285
rect 2273 283 2276 295
rect 2232 282 2261 283
rect 2256 279 2261 282
rect 2273 279 2279 283
rect 2256 278 2259 279
rect 2222 274 2232 278
rect 2246 274 2259 278
rect 2273 275 2276 279
rect 2220 257 2224 267
rect 2246 268 2250 274
rect 2266 257 2269 271
rect 2289 270 2292 334
rect 2329 327 2332 388
rect 2329 324 2398 327
rect 2340 318 2344 324
rect 2383 318 2386 324
rect 2333 299 2335 303
rect 2363 300 2367 309
rect 2391 302 2394 314
rect 2374 300 2379 302
rect 2361 298 2379 300
rect 2391 298 2396 302
rect 2361 296 2377 298
rect 2334 292 2354 295
rect 2361 289 2364 296
rect 2391 294 2394 298
rect 2352 286 2364 289
rect 2352 285 2356 286
rect 2384 285 2387 290
rect 2380 282 2387 285
rect 2340 270 2344 276
rect 2363 270 2367 276
rect 2380 270 2383 282
rect 2289 267 2376 270
rect 2289 257 2292 267
rect 2381 267 2383 270
rect 2220 254 2292 257
rect 2423 251 2430 577
rect 3174 544 3338 547
rect 2962 485 2973 489
rect 3174 489 3177 544
rect 3210 534 3214 544
rect 3240 534 3244 544
rect 3270 534 3274 544
rect 3295 534 3299 544
rect 3223 514 3227 530
rect 3255 514 3259 530
rect 3285 514 3289 530
rect 3311 514 3315 530
rect 3223 510 3302 514
rect 3311 510 3317 514
rect 3285 499 3289 510
rect 3311 505 3315 510
rect 2978 486 3177 489
rect 3210 489 3214 495
rect 3295 489 3299 495
rect 3335 495 3338 544
rect 3335 492 3724 495
rect 3210 486 3326 489
rect 2978 485 2987 486
rect 2968 480 2971 485
rect 2976 464 2979 476
rect 3210 474 3214 486
rect 3011 470 3214 474
rect 2976 460 2981 464
rect 2976 456 2979 460
rect 2969 447 2972 452
rect 3011 447 3014 470
rect 3233 469 3237 472
rect 3248 469 3252 472
rect 3263 469 3267 472
rect 3277 469 3281 472
rect 2968 444 2981 447
rect 2986 444 3014 447
rect 2964 419 2972 423
rect 2977 419 2989 423
rect 2970 414 2973 419
rect 2978 398 2981 410
rect 2978 394 2991 398
rect 2978 390 2981 394
rect 2971 381 2974 386
rect 3323 385 3326 486
rect 3335 447 3338 492
rect 3660 484 3664 492
rect 3720 484 3724 492
rect 3712 465 3716 480
rect 3733 469 3737 480
rect 3733 465 3742 469
rect 3673 461 3726 465
rect 3673 457 3677 461
rect 3699 457 3703 461
rect 3733 457 3737 465
rect 3335 444 3456 447
rect 3341 434 3345 444
rect 3374 434 3378 444
rect 3403 434 3407 444
rect 3412 434 3416 444
rect 3356 414 3361 430
rect 3389 414 3393 430
rect 3428 414 3432 430
rect 3356 410 3419 414
rect 3428 410 3434 414
rect 3403 399 3407 410
rect 3428 405 3432 410
rect 3453 409 3456 444
rect 3660 445 3664 450
rect 3686 445 3690 450
rect 3712 445 3716 453
rect 3720 445 3724 453
rect 3660 442 3724 445
rect 3453 406 3586 409
rect 3341 385 3345 395
rect 3412 385 3416 395
rect 3479 396 3483 406
rect 3512 396 3516 406
rect 3538 396 3542 406
rect 3323 382 3453 385
rect 2970 378 2981 381
rect 2967 352 2972 356
rect 2977 352 2992 356
rect 3384 359 3388 372
rect 3252 356 3388 359
rect 2973 347 2976 352
rect 3394 352 3398 371
rect 3267 349 3398 352
rect 3450 347 3453 382
rect 3494 376 3499 392
rect 3529 376 3533 392
rect 3554 376 3558 392
rect 3494 372 3545 376
rect 3554 372 3560 376
rect 3529 361 3533 372
rect 3554 367 3558 372
rect 3583 366 3586 406
rect 3583 362 3675 366
rect 3479 347 3483 357
rect 3538 347 3542 357
rect 3608 356 3612 362
rect 3450 344 3576 347
rect 2981 331 2984 343
rect 3043 334 3487 338
rect 3043 331 3047 334
rect 2981 327 3047 331
rect 2206 247 2207 251
rect 2211 247 2430 251
rect 2206 243 2430 247
rect 2981 323 2984 327
rect 2443 184 2447 322
rect 3522 325 3526 333
rect 3253 322 3526 325
rect 3573 319 3576 344
rect 3619 336 3623 353
rect 3629 356 3633 362
rect 3656 357 3659 362
rect 3640 336 3644 353
rect 3664 341 3667 353
rect 3647 337 3652 341
rect 3664 337 3668 341
rect 3647 336 3650 337
rect 3619 332 3650 336
rect 3664 333 3667 337
rect 3608 319 3612 325
rect 3640 326 3644 332
rect 3657 319 3660 329
rect 3717 319 3720 442
rect 2974 314 2977 319
rect 3573 316 3720 319
rect 2973 311 2981 314
rect 2967 285 2972 289
rect 2977 285 2992 289
rect 2973 280 2976 285
rect 2981 264 2984 276
rect 2981 260 3424 264
rect 2981 256 2984 260
rect 2974 247 2977 252
rect 2973 244 2981 247
rect 2443 180 2972 184
rect 2180 127 2276 130
rect 2091 119 2131 123
rect 2091 95 2095 119
rect 2091 78 2095 91
rect 2069 75 2095 78
rect 2069 67 2072 75
rect 2069 3 2072 62
rect 2091 64 2095 75
rect 2100 112 2118 116
rect 2100 95 2104 112
rect 2119 95 2123 111
rect 2100 64 2104 91
rect 2110 64 2114 91
rect 2119 64 2123 91
rect 2127 79 2131 119
rect 2180 111 2183 127
rect 2135 107 2183 111
rect 2135 95 2139 107
rect 2154 95 2158 107
rect 2127 75 2137 79
rect 2144 71 2148 91
rect 2127 67 2148 71
rect 2110 57 2114 60
rect 2127 57 2131 67
rect 2144 64 2148 67
rect 2163 79 2167 91
rect 2163 75 2166 79
rect 2163 64 2167 75
rect 2110 53 2131 57
rect 2135 57 2139 60
rect 2154 57 2158 60
rect 2135 53 2153 57
rect 2075 46 2115 49
rect 2075 37 2078 46
rect 2180 33 2183 107
rect 2228 115 2268 119
rect 2228 91 2232 115
rect 2228 74 2232 87
rect 2214 71 2232 74
rect 2228 60 2232 71
rect 2237 108 2260 112
rect 2237 91 2241 108
rect 2256 91 2260 108
rect 2237 60 2241 87
rect 2247 60 2251 87
rect 2256 60 2260 87
rect 2264 75 2268 115
rect 2272 107 2276 127
rect 2272 103 2335 107
rect 2272 91 2276 103
rect 2291 91 2295 103
rect 2264 71 2274 75
rect 2281 67 2285 87
rect 2264 63 2285 67
rect 2247 53 2251 56
rect 2264 53 2268 63
rect 2281 60 2285 63
rect 2300 75 2304 87
rect 2300 71 2303 75
rect 2300 60 2304 71
rect 2247 49 2268 53
rect 2272 53 2276 56
rect 2291 53 2295 56
rect 2272 49 2295 53
rect 2214 42 2250 45
rect 2272 39 2275 49
rect 2191 36 2275 39
rect 2075 12 2078 32
rect 2115 29 2200 33
rect 2121 23 2125 29
rect 2075 8 2125 12
rect 2133 10 2137 20
rect 2147 23 2151 29
rect 2166 24 2169 29
rect 2197 23 2200 29
rect 2133 8 2160 10
rect 2174 8 2177 20
rect 2197 19 2287 23
rect 2223 13 2227 19
rect 2133 7 2162 8
rect 2157 4 2162 7
rect 2174 4 2193 8
rect 2157 3 2160 4
rect 2069 -1 2133 3
rect 2147 -1 2160 3
rect 2174 0 2177 4
rect 2121 -16 2125 -8
rect 2147 -7 2151 -1
rect 2167 -15 2170 -4
rect 2125 -20 2167 -18
rect 2125 -21 2170 -20
rect 2190 -26 2193 4
rect 2210 2 2214 10
rect 2214 -2 2227 2
rect 2235 0 2239 10
rect 2249 13 2253 19
rect 2268 14 2271 19
rect 2235 -2 2262 0
rect 2276 -2 2279 10
rect 2235 -3 2264 -2
rect 2259 -6 2264 -3
rect 2276 -6 2282 -2
rect 2259 -7 2262 -6
rect 2225 -11 2235 -7
rect 2249 -11 2262 -7
rect 2276 -10 2279 -6
rect 2223 -28 2227 -18
rect 2249 -17 2253 -11
rect 2269 -28 2272 -14
rect 2292 -15 2295 49
rect 2332 42 2335 103
rect 2443 42 2447 180
rect 2891 162 2931 166
rect 2891 138 2895 162
rect 2891 121 2895 134
rect 2878 118 2895 121
rect 2891 107 2895 118
rect 2900 155 2919 159
rect 2900 138 2904 155
rect 2919 138 2923 154
rect 2900 107 2904 134
rect 2910 107 2914 134
rect 2919 107 2923 134
rect 2927 122 2931 162
rect 2954 154 2958 180
rect 2977 180 3010 184
rect 2991 175 2994 180
rect 2999 159 3002 171
rect 2985 155 2987 159
rect 2999 155 3109 159
rect 2935 150 2958 154
rect 2999 151 3002 155
rect 2935 138 2939 150
rect 2954 138 2958 150
rect 2992 142 2995 147
rect 2980 139 2995 142
rect 2927 118 2937 122
rect 2944 114 2948 134
rect 2927 110 2948 114
rect 2910 100 2914 103
rect 2927 100 2931 110
rect 2944 107 2948 110
rect 2963 122 2967 134
rect 2963 118 2966 122
rect 2963 107 2967 118
rect 2910 96 2931 100
rect 2935 100 2939 103
rect 2954 100 2958 103
rect 2980 101 2985 139
rect 2980 100 2981 101
rect 2935 96 2981 100
rect 2877 89 2915 92
rect 2877 79 2880 89
rect 2332 39 2447 42
rect 2823 76 2880 79
rect 2343 33 2347 39
rect 2386 33 2389 39
rect 2336 14 2338 18
rect 2366 15 2370 24
rect 2394 17 2397 29
rect 2377 15 2382 17
rect 2364 13 2382 15
rect 2394 13 2419 17
rect 2364 11 2380 13
rect 2337 7 2357 10
rect 2364 4 2367 11
rect 2394 9 2397 13
rect 2355 1 2367 4
rect 2355 0 2359 1
rect 2387 0 2390 5
rect 2383 -3 2390 0
rect 2343 -15 2347 -9
rect 2366 -15 2370 -9
rect 2383 -15 2386 -3
rect 2292 -18 2376 -15
rect 2292 -28 2295 -18
rect 2381 -18 2386 -15
rect 2223 -31 2295 -28
rect 2009 -72 2029 -71
rect 1212 -73 1241 -72
rect 1236 -76 1241 -73
rect 1253 -76 2029 -72
rect 1236 -77 1239 -76
rect 1202 -81 1212 -77
rect 1226 -81 1239 -77
rect 1253 -80 1256 -76
rect 1200 -98 1204 -88
rect 1226 -87 1230 -81
rect 1246 -98 1249 -84
rect 1200 -101 1238 -98
rect 1243 -101 1249 -98
rect 487 -134 1792 -131
rect 417 -138 422 -134
rect 434 -138 455 -134
rect 417 -139 420 -138
rect 383 -143 420 -139
rect 434 -142 437 -138
rect 372 -163 376 -150
rect 383 -156 387 -150
rect 398 -156 402 -150
rect 409 -149 413 -143
rect 427 -151 430 -146
rect 383 -160 402 -156
rect 423 -154 453 -151
rect 423 -163 426 -154
rect 372 -166 426 -163
rect 69 -170 101 -166
rect 113 -170 183 -166
rect 75 -267 82 -170
rect 113 -174 116 -170
rect 106 -181 109 -178
rect 369 -181 439 -178
rect 86 -201 92 -188
rect 372 -188 376 -181
rect 86 -205 189 -201
rect 195 -205 376 -201
rect 383 -208 387 -191
rect 398 -188 402 -181
rect 420 -182 439 -181
rect 426 -187 429 -182
rect 444 -182 445 -178
rect 400 -205 402 -201
rect 409 -208 413 -191
rect 417 -207 422 -203
rect 417 -208 420 -207
rect 383 -212 420 -208
rect 434 -211 437 -191
rect 372 -232 376 -219
rect 383 -225 387 -219
rect 398 -225 402 -219
rect 409 -218 413 -212
rect 427 -220 430 -215
rect 449 -220 452 -154
rect 487 -178 491 -134
rect 537 -140 541 -134
rect 580 -140 583 -134
rect 685 -135 1792 -134
rect 685 -141 689 -135
rect 531 -159 532 -155
rect 560 -158 564 -149
rect 588 -156 591 -144
rect 697 -154 701 -144
rect 711 -141 715 -135
rect 730 -140 733 -135
rect 823 -141 827 -135
rect 697 -156 724 -154
rect 738 -156 741 -144
rect 835 -154 839 -144
rect 849 -141 853 -135
rect 868 -140 871 -135
rect 969 -141 973 -135
rect 571 -158 576 -156
rect 558 -160 576 -158
rect 588 -160 593 -156
rect 697 -157 726 -156
rect 721 -160 726 -157
rect 738 -160 744 -156
rect 835 -156 862 -154
rect 876 -156 879 -144
rect 981 -154 985 -144
rect 995 -141 999 -135
rect 1014 -140 1017 -135
rect 1093 -141 1097 -135
rect 835 -157 864 -156
rect 859 -160 864 -157
rect 876 -160 882 -156
rect 558 -162 574 -160
rect 509 -166 517 -163
rect 521 -166 551 -163
rect 558 -169 561 -162
rect 588 -164 591 -160
rect 721 -161 724 -160
rect 688 -165 697 -161
rect 711 -165 724 -161
rect 738 -164 741 -160
rect 549 -172 561 -169
rect 549 -173 553 -172
rect 581 -173 584 -168
rect 577 -176 584 -173
rect 383 -229 402 -225
rect 423 -223 449 -220
rect 423 -232 426 -223
rect 372 -235 426 -232
rect 366 -247 441 -244
rect 372 -254 376 -247
rect 75 -271 376 -267
rect 343 -333 350 -271
rect 383 -274 387 -257
rect 398 -254 402 -247
rect 420 -248 441 -247
rect 426 -253 429 -248
rect 400 -271 402 -267
rect 409 -274 413 -257
rect 434 -269 437 -257
rect 417 -273 422 -269
rect 434 -273 438 -269
rect 417 -274 420 -273
rect 383 -278 420 -274
rect 434 -277 437 -273
rect 372 -299 376 -285
rect 383 -291 387 -285
rect 398 -291 402 -285
rect 409 -284 413 -278
rect 427 -286 430 -281
rect 449 -286 452 -225
rect 487 -244 491 -183
rect 537 -188 541 -182
rect 560 -188 564 -182
rect 577 -182 580 -176
rect 685 -182 689 -172
rect 711 -171 715 -165
rect 859 -161 862 -160
rect 826 -165 835 -161
rect 849 -165 862 -161
rect 876 -164 879 -160
rect 981 -156 1008 -154
rect 1022 -156 1025 -144
rect 1105 -154 1109 -144
rect 1119 -141 1123 -135
rect 1138 -140 1141 -135
rect 1318 -141 1322 -135
rect 1105 -156 1132 -154
rect 1146 -156 1149 -144
rect 1330 -154 1334 -144
rect 1344 -141 1348 -135
rect 1363 -140 1366 -135
rect 1465 -141 1469 -135
rect 1330 -156 1357 -154
rect 981 -157 1010 -156
rect 1005 -160 1010 -157
rect 1022 -160 1028 -156
rect 731 -182 734 -168
rect 823 -182 827 -172
rect 849 -171 853 -165
rect 1005 -161 1008 -160
rect 971 -165 981 -161
rect 995 -165 1008 -161
rect 1022 -164 1025 -160
rect 1105 -157 1134 -156
rect 1129 -160 1134 -157
rect 1146 -160 1152 -156
rect 869 -182 872 -168
rect 969 -182 973 -172
rect 995 -171 999 -165
rect 1129 -161 1132 -160
rect 1095 -165 1105 -161
rect 1119 -165 1132 -161
rect 1146 -164 1149 -160
rect 1330 -157 1359 -156
rect 1354 -160 1359 -157
rect 1015 -182 1018 -168
rect 1093 -182 1097 -172
rect 1119 -171 1123 -165
rect 1354 -161 1357 -160
rect 1320 -165 1330 -161
rect 1344 -165 1357 -161
rect 1371 -164 1374 -144
rect 1477 -154 1481 -144
rect 1491 -141 1495 -135
rect 1510 -140 1513 -135
rect 1604 -141 1608 -135
rect 1477 -156 1504 -154
rect 1518 -156 1521 -144
rect 1616 -154 1620 -144
rect 1630 -141 1634 -135
rect 1649 -140 1652 -135
rect 1728 -141 1732 -135
rect 1477 -157 1506 -156
rect 1501 -160 1506 -157
rect 1518 -160 1524 -156
rect 1616 -156 1643 -154
rect 1657 -156 1660 -144
rect 1740 -154 1744 -144
rect 1754 -141 1758 -135
rect 1773 -140 1776 -135
rect 1616 -157 1645 -156
rect 1640 -160 1645 -157
rect 1657 -160 1663 -156
rect 1740 -156 1767 -154
rect 1781 -156 1784 -144
rect 1740 -157 1769 -156
rect 1764 -160 1769 -157
rect 1781 -160 1787 -156
rect 1139 -182 1142 -168
rect 1318 -182 1322 -172
rect 1344 -171 1348 -165
rect 1501 -161 1504 -160
rect 1467 -165 1477 -161
rect 1491 -165 1504 -161
rect 1518 -164 1521 -160
rect 1364 -182 1367 -168
rect 1465 -182 1469 -172
rect 1491 -171 1495 -165
rect 1640 -161 1643 -160
rect 1606 -165 1616 -161
rect 1630 -165 1643 -161
rect 1657 -164 1660 -160
rect 1511 -182 1514 -168
rect 1604 -182 1608 -172
rect 1630 -171 1634 -165
rect 1764 -161 1767 -160
rect 1730 -165 1740 -161
rect 1754 -165 1767 -161
rect 1781 -164 1784 -160
rect 1650 -182 1653 -168
rect 1728 -182 1732 -172
rect 1754 -171 1758 -165
rect 1774 -182 1777 -168
rect 577 -185 1238 -182
rect 577 -188 580 -185
rect 1243 -185 1852 -182
rect 539 -191 580 -188
rect 490 -249 491 -244
rect 383 -295 402 -291
rect 423 -289 452 -286
rect 423 -299 426 -289
rect 372 -302 426 -299
rect 366 -313 440 -310
rect 372 -320 376 -313
rect 343 -337 376 -333
rect 383 -340 387 -323
rect 398 -320 402 -313
rect 420 -314 440 -313
rect 426 -319 429 -314
rect 400 -337 402 -333
rect 409 -340 413 -323
rect 434 -335 437 -323
rect 417 -339 422 -335
rect 434 -339 439 -335
rect 417 -340 420 -339
rect 383 -344 420 -340
rect 434 -343 437 -339
rect 372 -367 376 -351
rect 383 -357 387 -351
rect 398 -357 402 -351
rect 409 -350 413 -344
rect 427 -352 430 -347
rect 449 -352 452 -289
rect 487 -264 491 -249
rect 487 -267 1787 -264
rect 487 -310 491 -267
rect 680 -268 1787 -267
rect 680 -274 684 -268
rect 692 -287 696 -277
rect 706 -274 710 -268
rect 725 -273 728 -268
rect 818 -274 822 -268
rect 692 -289 719 -287
rect 733 -289 736 -277
rect 830 -287 834 -277
rect 844 -274 848 -268
rect 863 -273 866 -268
rect 964 -274 968 -268
rect 830 -289 857 -287
rect 871 -289 874 -277
rect 976 -287 980 -277
rect 990 -274 994 -268
rect 1009 -273 1012 -268
rect 1088 -274 1092 -268
rect 976 -289 1003 -287
rect 1017 -289 1020 -277
rect 1100 -287 1104 -277
rect 1114 -274 1118 -268
rect 1133 -273 1136 -268
rect 1313 -274 1317 -268
rect 1100 -289 1127 -287
rect 1141 -289 1144 -277
rect 1325 -287 1329 -277
rect 1339 -274 1343 -268
rect 1358 -273 1361 -268
rect 1460 -274 1464 -268
rect 1325 -289 1352 -287
rect 1366 -289 1369 -277
rect 1472 -287 1476 -277
rect 1486 -274 1490 -268
rect 1505 -273 1508 -268
rect 1599 -274 1603 -268
rect 1472 -289 1499 -287
rect 1513 -289 1516 -277
rect 1611 -287 1615 -277
rect 1625 -274 1629 -268
rect 1644 -273 1647 -268
rect 1723 -274 1727 -268
rect 1611 -289 1638 -287
rect 1652 -289 1655 -277
rect 1735 -287 1739 -277
rect 1749 -274 1753 -268
rect 1768 -273 1771 -268
rect 1735 -289 1762 -287
rect 1776 -289 1779 -277
rect 2823 -289 2826 76
rect 2956 19 2972 23
rect 2893 1 2933 5
rect 2893 -23 2897 1
rect 2893 -40 2897 -27
rect 2880 -43 2897 -40
rect 2893 -54 2897 -43
rect 2902 -6 2921 -2
rect 2902 -23 2906 -6
rect 2921 -23 2925 -7
rect 2902 -54 2906 -27
rect 2912 -54 2916 -27
rect 2921 -54 2925 -27
rect 2929 -39 2933 1
rect 2956 -7 2960 19
rect 2977 19 3007 23
rect 2993 14 2996 19
rect 3001 -2 3004 10
rect 2987 -6 2989 -2
rect 3001 -4 3071 -2
rect 2937 -11 2960 -7
rect 3001 -7 3072 -4
rect 3001 -10 3004 -7
rect 2937 -23 2941 -11
rect 2956 -23 2960 -11
rect 2994 -19 2997 -14
rect 2929 -43 2939 -39
rect 2946 -47 2950 -27
rect 2929 -51 2950 -47
rect 2912 -61 2916 -58
rect 2929 -61 2933 -51
rect 2946 -54 2950 -51
rect 2965 -39 2969 -27
rect 2987 -22 2997 -19
rect 2965 -43 2968 -39
rect 2965 -54 2969 -43
rect 2912 -65 2933 -61
rect 2937 -61 2941 -58
rect 2956 -61 2960 -58
rect 2982 -61 2987 -24
rect 2937 -65 2987 -61
rect 2879 -72 2917 -69
rect 2879 -79 2882 -72
rect 3063 -73 3072 -7
rect 3100 -53 3109 155
rect 3502 48 3506 312
rect 3634 300 3638 307
rect 3154 45 3506 48
rect 3585 -30 3691 -27
rect 3588 -40 3592 -30
rect 3621 -40 3625 -30
rect 3650 -40 3654 -30
rect 3659 -40 3663 -30
rect 3688 -32 3691 -30
rect 3688 -36 3781 -32
rect 3100 -58 3247 -53
rect 3252 -58 3546 -53
rect 3101 -59 3546 -58
rect 692 -290 721 -289
rect 716 -293 721 -290
rect 733 -293 745 -289
rect 830 -290 859 -289
rect 854 -293 859 -290
rect 871 -293 884 -289
rect 976 -290 1005 -289
rect 1000 -293 1005 -290
rect 1017 -293 1027 -289
rect 1100 -290 1129 -289
rect 1124 -293 1129 -290
rect 1141 -293 1151 -289
rect 1325 -290 1354 -289
rect 1349 -293 1354 -290
rect 1366 -293 1378 -289
rect 1472 -290 1501 -289
rect 1496 -293 1501 -290
rect 1513 -293 1527 -289
rect 1611 -290 1640 -289
rect 1635 -293 1640 -290
rect 1652 -291 1668 -289
rect 1735 -290 1764 -289
rect 1652 -293 1664 -291
rect 716 -294 719 -293
rect 683 -298 692 -294
rect 706 -298 719 -294
rect 733 -297 736 -293
rect 490 -315 491 -310
rect 680 -314 684 -305
rect 706 -304 710 -298
rect 854 -294 857 -293
rect 821 -298 830 -294
rect 844 -298 857 -294
rect 871 -297 874 -293
rect 383 -361 402 -357
rect 423 -355 452 -352
rect 423 -367 426 -355
rect 372 -370 426 -367
rect 71 -403 105 -402
rect 394 -402 399 -370
rect 487 -373 491 -315
rect 599 -315 684 -314
rect 726 -315 729 -301
rect 818 -315 822 -305
rect 844 -304 848 -298
rect 1000 -294 1003 -293
rect 965 -298 976 -294
rect 990 -298 1003 -294
rect 1017 -297 1020 -293
rect 864 -315 867 -301
rect 964 -315 968 -305
rect 990 -304 994 -298
rect 1124 -294 1127 -293
rect 1089 -298 1100 -294
rect 1114 -298 1127 -294
rect 1141 -297 1144 -293
rect 1010 -315 1013 -301
rect 1088 -315 1092 -305
rect 1114 -304 1118 -298
rect 1349 -294 1352 -293
rect 1314 -298 1325 -294
rect 1339 -298 1352 -294
rect 1366 -297 1369 -293
rect 1134 -315 1137 -301
rect 1313 -315 1317 -305
rect 1339 -304 1343 -298
rect 1496 -294 1499 -293
rect 1462 -298 1472 -294
rect 1486 -298 1499 -294
rect 1513 -297 1516 -293
rect 1359 -315 1362 -301
rect 1460 -315 1464 -305
rect 1486 -304 1490 -298
rect 1635 -294 1638 -293
rect 1601 -298 1611 -294
rect 1625 -298 1638 -294
rect 1652 -297 1655 -293
rect 1759 -293 1764 -290
rect 1776 -293 2826 -289
rect 1506 -315 1509 -301
rect 1599 -315 1603 -305
rect 1625 -304 1629 -298
rect 1759 -294 1762 -293
rect 1725 -298 1735 -294
rect 1749 -298 1762 -294
rect 1776 -297 1779 -293
rect 1645 -315 1648 -301
rect 1723 -315 1727 -305
rect 1749 -304 1753 -298
rect 1769 -315 1772 -301
rect 599 -318 1772 -315
rect 2739 -350 2762 -346
rect 487 -378 635 -373
rect 110 -403 466 -402
rect 71 -405 466 -403
rect 462 -454 466 -405
rect 631 -403 635 -378
rect 2773 -378 2777 -375
rect 631 -406 1809 -403
rect 676 -407 1809 -406
rect 676 -413 680 -407
rect 688 -426 692 -416
rect 702 -413 706 -407
rect 721 -412 724 -407
rect 814 -413 818 -407
rect 688 -428 715 -426
rect 729 -428 732 -416
rect 826 -426 830 -416
rect 840 -413 844 -407
rect 859 -412 862 -407
rect 960 -413 964 -407
rect 826 -428 853 -426
rect 867 -428 870 -416
rect 972 -426 976 -416
rect 986 -413 990 -407
rect 1005 -412 1008 -407
rect 1084 -413 1088 -407
rect 972 -428 999 -426
rect 1013 -428 1016 -416
rect 1096 -426 1100 -416
rect 1110 -413 1114 -407
rect 1129 -412 1132 -407
rect 1309 -413 1313 -407
rect 688 -429 717 -428
rect 712 -432 717 -429
rect 729 -432 734 -428
rect 826 -429 855 -428
rect 850 -432 855 -429
rect 867 -432 873 -428
rect 712 -433 715 -432
rect 678 -437 688 -433
rect 702 -437 715 -433
rect 729 -436 732 -432
rect 676 -454 680 -444
rect 702 -443 706 -437
rect 850 -433 853 -432
rect 816 -437 826 -433
rect 840 -437 853 -433
rect 867 -436 870 -432
rect 972 -429 1001 -428
rect 996 -432 1001 -429
rect 1013 -432 1019 -428
rect 1096 -428 1123 -426
rect 1137 -428 1140 -416
rect 1321 -426 1325 -416
rect 1335 -413 1339 -407
rect 1354 -412 1357 -407
rect 1456 -413 1460 -407
rect 1321 -428 1348 -426
rect 1362 -428 1365 -416
rect 1468 -426 1472 -416
rect 1482 -413 1486 -407
rect 1501 -412 1504 -407
rect 1595 -413 1599 -407
rect 1468 -428 1495 -426
rect 1509 -428 1512 -416
rect 1607 -426 1611 -416
rect 1621 -413 1625 -407
rect 1640 -412 1643 -407
rect 1719 -413 1723 -407
rect 1607 -428 1634 -426
rect 1648 -428 1651 -416
rect 1731 -426 1735 -416
rect 1745 -413 1749 -407
rect 1764 -412 1767 -407
rect 1731 -428 1758 -426
rect 1772 -428 1775 -416
rect 1096 -429 1125 -428
rect 1120 -432 1125 -429
rect 1137 -432 1143 -428
rect 722 -454 725 -440
rect 814 -454 818 -444
rect 840 -443 844 -437
rect 996 -433 999 -432
rect 961 -437 972 -433
rect 986 -437 999 -433
rect 1013 -436 1016 -432
rect 860 -454 863 -440
rect 960 -454 964 -444
rect 986 -443 990 -437
rect 1120 -433 1123 -432
rect 1085 -437 1096 -433
rect 1110 -437 1123 -433
rect 1137 -436 1140 -432
rect 1321 -429 1350 -428
rect 1345 -432 1350 -429
rect 1362 -432 1367 -428
rect 1468 -429 1497 -428
rect 1492 -432 1497 -429
rect 1509 -432 1514 -428
rect 1607 -429 1636 -428
rect 1631 -432 1636 -429
rect 1648 -432 1653 -428
rect 1731 -429 1760 -428
rect 1755 -432 1760 -429
rect 1772 -432 1777 -428
rect 1006 -454 1009 -440
rect 1084 -454 1088 -444
rect 1110 -443 1114 -437
rect 1345 -433 1348 -432
rect 1310 -437 1321 -433
rect 1335 -437 1348 -433
rect 1362 -436 1365 -432
rect 1130 -454 1133 -440
rect 1309 -454 1313 -444
rect 1335 -443 1339 -437
rect 1492 -433 1495 -432
rect 1458 -437 1468 -433
rect 1482 -437 1495 -433
rect 1509 -436 1512 -432
rect 1355 -454 1358 -440
rect 1456 -454 1460 -444
rect 1482 -443 1486 -437
rect 1631 -433 1634 -432
rect 1597 -437 1607 -433
rect 1621 -437 1634 -433
rect 1648 -436 1651 -432
rect 1502 -454 1505 -440
rect 1595 -454 1599 -444
rect 1621 -443 1625 -437
rect 1755 -433 1758 -432
rect 1721 -437 1731 -433
rect 1745 -437 1758 -433
rect 1772 -436 1775 -432
rect 1641 -454 1644 -440
rect 1719 -454 1723 -444
rect 1745 -443 1749 -437
rect 1765 -454 1768 -440
rect 1806 -447 1809 -407
rect 2728 -442 2797 -439
rect 1806 -451 1909 -447
rect 462 -457 1768 -454
rect 1765 -498 1768 -457
rect 1835 -457 1839 -451
rect 1847 -470 1851 -460
rect 1861 -457 1865 -451
rect 1880 -456 1883 -451
rect 1847 -472 1874 -470
rect 1888 -472 1891 -460
rect 1847 -473 1876 -472
rect 1871 -476 1876 -473
rect 1888 -476 1895 -472
rect 1871 -477 1874 -476
rect 1838 -481 1847 -477
rect 1861 -481 1874 -477
rect 1888 -480 1891 -476
rect 1835 -498 1839 -488
rect 1861 -487 1865 -481
rect 1881 -498 1884 -484
rect 1765 -501 1884 -498
rect 1765 -603 1768 -501
rect 1906 -552 1909 -451
rect 2752 -535 2756 -533
rect 1829 -556 1909 -552
rect 1835 -562 1839 -556
rect 1847 -575 1851 -565
rect 1861 -562 1865 -556
rect 1880 -561 1883 -556
rect 1847 -577 1874 -575
rect 1888 -577 1891 -565
rect 1847 -578 1876 -577
rect 1871 -581 1876 -578
rect 1888 -581 1895 -577
rect 1871 -582 1874 -581
rect 1839 -586 1847 -582
rect 1861 -586 1874 -582
rect 1888 -585 1891 -581
rect 1835 -603 1839 -593
rect 1861 -592 1865 -586
rect 1881 -603 1884 -589
rect 1765 -606 1884 -603
rect 1765 -725 1768 -606
rect 1906 -674 1909 -556
rect 2823 -668 2826 -293
rect 2841 -82 2882 -79
rect 3063 -78 3262 -73
rect 3267 -78 3525 -73
rect 3063 -80 3525 -78
rect 3063 -81 3072 -80
rect 2841 -525 2844 -82
rect 3522 -102 3525 -80
rect 3543 -95 3546 -59
rect 3603 -60 3608 -44
rect 3636 -60 3640 -44
rect 3675 -60 3679 -44
rect 3703 -42 3707 -36
rect 3696 -59 3707 -55
rect 3696 -60 3699 -59
rect 3603 -64 3666 -60
rect 3675 -64 3699 -60
rect 3714 -62 3718 -45
rect 3729 -42 3733 -36
rect 3762 -41 3765 -36
rect 3729 -59 3733 -55
rect 3740 -62 3744 -45
rect 3770 -57 3773 -45
rect 3753 -61 3758 -57
rect 3770 -61 3777 -57
rect 3753 -62 3756 -61
rect 3650 -75 3654 -64
rect 3675 -69 3679 -64
rect 3714 -66 3756 -62
rect 3770 -65 3773 -61
rect 3588 -89 3592 -79
rect 3659 -86 3663 -79
rect 3703 -86 3707 -73
rect 3740 -72 3744 -66
rect 3659 -87 3707 -86
rect 3763 -87 3766 -69
rect 3659 -89 3766 -87
rect 3588 -92 3658 -89
rect 3663 -90 3766 -89
rect 3543 -98 3570 -95
rect 3522 -105 3570 -102
rect 3424 -113 3570 -110
rect 2897 -121 2908 -117
rect 2955 -135 2972 -131
rect 2892 -153 2932 -149
rect 2892 -177 2896 -153
rect 2892 -194 2896 -181
rect 2879 -197 2896 -194
rect 2892 -208 2896 -197
rect 2901 -160 2920 -156
rect 2901 -177 2905 -160
rect 2920 -177 2924 -161
rect 2901 -208 2905 -181
rect 2911 -208 2915 -181
rect 2920 -208 2924 -181
rect 2928 -193 2932 -153
rect 2955 -161 2959 -135
rect 2977 -135 3011 -131
rect 2992 -140 2995 -135
rect 3000 -156 3003 -144
rect 2986 -160 2988 -156
rect 3000 -160 3276 -156
rect 3424 -156 3427 -113
rect 3281 -160 3427 -156
rect 3496 -122 3570 -119
rect 2936 -165 2959 -161
rect 3000 -164 3003 -160
rect 2936 -177 2940 -165
rect 2955 -177 2959 -165
rect 2993 -173 2996 -168
rect 2928 -197 2938 -193
rect 2945 -201 2949 -181
rect 2928 -205 2949 -201
rect 2911 -215 2915 -212
rect 2928 -215 2932 -205
rect 2945 -208 2949 -205
rect 2964 -193 2968 -181
rect 2986 -176 2996 -173
rect 2964 -197 2967 -193
rect 2964 -208 2968 -197
rect 2911 -219 2932 -215
rect 2936 -215 2940 -212
rect 2955 -215 2959 -212
rect 2981 -215 2986 -178
rect 2936 -219 2986 -215
rect 2878 -226 2916 -223
rect 2878 -234 2881 -226
rect 2852 -237 2881 -234
rect 2852 -385 2855 -237
rect 2955 -283 2972 -279
rect 2892 -301 2932 -297
rect 2892 -325 2896 -301
rect 2892 -342 2896 -329
rect 2879 -345 2896 -342
rect 2892 -356 2896 -345
rect 2901 -308 2920 -304
rect 2901 -325 2905 -308
rect 2920 -325 2924 -309
rect 2901 -356 2905 -329
rect 2911 -356 2915 -329
rect 2920 -356 2924 -329
rect 2928 -341 2932 -301
rect 2955 -309 2959 -283
rect 2977 -283 3011 -279
rect 2992 -288 2995 -283
rect 3000 -304 3003 -292
rect 3496 -304 3502 -122
rect 2986 -308 2988 -304
rect 3000 -308 3502 -304
rect 3592 -288 3715 -285
rect 2936 -313 2959 -309
rect 3000 -312 3003 -308
rect 2936 -325 2940 -313
rect 2955 -325 2959 -313
rect 2993 -321 2996 -316
rect 2928 -345 2938 -341
rect 2945 -349 2949 -329
rect 2928 -353 2949 -349
rect 2911 -363 2915 -360
rect 2928 -363 2932 -353
rect 2945 -356 2949 -353
rect 2964 -341 2968 -329
rect 2986 -324 2996 -321
rect 2964 -345 2967 -341
rect 2964 -356 2968 -345
rect 2911 -367 2932 -363
rect 2936 -363 2940 -360
rect 2955 -363 2959 -360
rect 2981 -363 2986 -326
rect 3592 -342 3595 -288
rect 3651 -296 3655 -288
rect 3711 -296 3715 -288
rect 3703 -315 3707 -300
rect 3724 -311 3728 -300
rect 3724 -315 3733 -311
rect 3664 -319 3717 -315
rect 3664 -323 3668 -319
rect 3690 -323 3694 -319
rect 3724 -323 3728 -315
rect 3651 -335 3655 -330
rect 3677 -335 3681 -330
rect 3703 -335 3707 -327
rect 3711 -335 3715 -327
rect 3651 -338 3715 -335
rect 3421 -345 3595 -342
rect 3425 -355 3429 -345
rect 3455 -355 3459 -345
rect 3485 -355 3489 -345
rect 3510 -355 3514 -345
rect 2936 -367 2986 -363
rect 2878 -374 2916 -371
rect 2878 -388 2881 -374
rect 3438 -375 3442 -359
rect 3470 -375 3474 -359
rect 3500 -375 3504 -359
rect 3526 -375 3530 -359
rect 3438 -379 3517 -375
rect 3526 -379 3532 -375
rect 2852 -461 2855 -389
rect 2878 -391 2907 -388
rect 2911 -391 3420 -388
rect 3500 -390 3504 -379
rect 3526 -384 3530 -379
rect 2962 -410 2972 -406
rect 2977 -410 2987 -406
rect 2968 -415 2971 -410
rect 2976 -431 2979 -419
rect 3387 -426 3390 -405
rect 3415 -421 3420 -391
rect 3425 -400 3429 -394
rect 3510 -400 3514 -394
rect 3664 -400 3667 -338
rect 3685 -353 3689 -347
rect 3425 -403 3667 -400
rect 3448 -421 3452 -418
rect 3415 -424 3452 -421
rect 3290 -429 3390 -426
rect 2932 -435 2951 -431
rect 2976 -435 3035 -431
rect 2976 -439 2979 -435
rect 3293 -439 3297 -429
rect 3326 -439 3330 -429
rect 3355 -439 3359 -429
rect 3364 -439 3368 -429
rect 2969 -448 2972 -443
rect 2968 -451 2981 -448
rect 3308 -459 3313 -443
rect 3341 -459 3345 -443
rect 3380 -459 3384 -443
rect 2852 -465 3275 -461
rect 3308 -463 3371 -459
rect 3380 -463 3386 -459
rect 2964 -476 2972 -472
rect 2977 -476 2989 -472
rect 2970 -481 2973 -476
rect 2978 -497 2981 -485
rect 2932 -501 2951 -497
rect 2978 -501 2992 -497
rect 2978 -505 2981 -501
rect 3149 -504 3233 -501
rect 2971 -514 2974 -509
rect 3152 -514 3156 -504
rect 3185 -514 3189 -504
rect 3211 -514 3215 -504
rect 3271 -505 3275 -465
rect 3355 -474 3359 -463
rect 3380 -468 3384 -463
rect 3293 -488 3297 -478
rect 3364 -488 3368 -478
rect 3455 -488 3458 -403
rect 3463 -426 3467 -418
rect 3293 -491 3458 -488
rect 3316 -505 3320 -501
rect 3271 -508 3320 -505
rect 3326 -513 3330 -491
rect 3336 -506 3340 -500
rect 3346 -506 3350 -500
rect 2970 -517 2981 -514
rect 2841 -528 2868 -525
rect 2874 -528 3140 -525
rect 2967 -543 2972 -539
rect 2977 -543 2992 -539
rect 2973 -548 2976 -543
rect 2850 -566 2856 -563
rect 2981 -564 2984 -552
rect 2924 -568 2951 -564
rect 2981 -568 2986 -564
rect 2981 -572 2984 -568
rect 2974 -581 2977 -576
rect 2973 -584 2981 -581
rect 3036 -582 3120 -578
rect 2967 -610 2972 -606
rect 3036 -606 3039 -582
rect 3057 -588 3061 -582
rect 2977 -610 3039 -606
rect 3068 -608 3072 -591
rect 3078 -588 3082 -582
rect 3105 -587 3108 -582
rect 3137 -582 3140 -528
rect 3167 -534 3172 -518
rect 3202 -534 3206 -518
rect 3227 -534 3231 -518
rect 3281 -516 3330 -513
rect 3167 -538 3218 -534
rect 3227 -538 3234 -534
rect 3202 -549 3206 -538
rect 3227 -543 3231 -538
rect 3152 -563 3156 -553
rect 3211 -563 3215 -553
rect 3281 -563 3284 -516
rect 3321 -527 3324 -525
rect 3478 -527 3482 -417
rect 3492 -425 3496 -417
rect 3321 -530 3482 -527
rect 3152 -566 3284 -563
rect 3175 -582 3179 -576
rect 3137 -585 3179 -582
rect 3089 -608 3093 -591
rect 3113 -603 3116 -591
rect 3096 -607 3101 -603
rect 3113 -607 3117 -603
rect 3096 -608 3099 -607
rect 2973 -615 2976 -610
rect 3068 -612 3099 -608
rect 3113 -611 3116 -607
rect 2981 -631 2984 -619
rect 3057 -626 3061 -619
rect 3089 -618 3093 -612
rect 3106 -626 3109 -615
rect 3186 -626 3189 -566
rect 3195 -581 3199 -577
rect 3057 -629 3189 -626
rect 2903 -635 2951 -631
rect 2981 -635 2987 -631
rect 2981 -639 2984 -635
rect 2974 -648 2977 -643
rect 3072 -648 3075 -629
rect 2973 -651 2981 -648
rect 2986 -651 3075 -648
rect 3083 -668 3087 -639
rect 2823 -671 3087 -668
rect 1829 -678 1909 -674
rect 1835 -684 1839 -678
rect 1847 -697 1851 -687
rect 1861 -684 1865 -678
rect 1880 -683 1883 -678
rect 1847 -699 1874 -697
rect 1888 -699 1891 -687
rect 1847 -700 1876 -699
rect 1871 -703 1876 -700
rect 1888 -703 1895 -699
rect 1871 -704 1874 -703
rect 1839 -708 1847 -704
rect 1861 -708 1874 -704
rect 1888 -707 1891 -703
rect 1835 -725 1839 -715
rect 1861 -714 1865 -708
rect 1881 -725 1884 -711
rect 1765 -728 1884 -725
rect 1765 -832 1768 -728
rect 1906 -781 1909 -678
rect 1829 -785 1909 -781
rect 1835 -791 1839 -785
rect 1847 -804 1851 -794
rect 1861 -791 1865 -785
rect 1880 -790 1883 -785
rect 1847 -806 1874 -804
rect 1888 -806 1891 -794
rect 1847 -807 1876 -806
rect 1871 -810 1876 -807
rect 1888 -810 1895 -806
rect 1871 -811 1874 -810
rect 1837 -815 1847 -811
rect 1861 -815 1874 -811
rect 1888 -814 1891 -810
rect 1835 -832 1839 -822
rect 1861 -821 1865 -815
rect 1881 -832 1884 -818
rect 3106 -832 3109 -629
rect 1765 -835 3109 -832
<< m2contact >>
rect 2120 951 2125 956
rect 2155 892 2160 897
rect 2067 876 2072 882
rect 2211 909 2216 914
rect 2211 882 2216 887
rect 2188 876 2193 881
rect 2211 850 2217 855
rect 2169 820 2174 825
rect 2284 834 2289 839
rect 2222 829 2227 834
rect 2190 809 2195 814
rect 2333 854 2338 859
rect 2334 845 2339 850
rect 2371 820 2376 825
rect 136 -74 141 -69
rect 366 -102 371 -97
rect 254 -116 260 -110
rect 86 -137 92 -131
rect 104 -132 109 -127
rect 121 -146 126 -141
rect 341 -144 347 -138
rect 394 -136 400 -129
rect 1456 50 1461 55
rect 1411 -16 1416 -11
rect 1604 47 1609 52
rect 1558 -18 1563 -13
rect 1756 47 1761 52
rect 1709 -19 1714 -14
rect 1908 46 1913 51
rect 1861 -20 1866 -15
rect 2118 675 2123 680
rect 2153 616 2158 621
rect 2067 597 2072 602
rect 2209 633 2214 638
rect 2209 606 2214 611
rect 2186 600 2191 605
rect 2209 574 2215 579
rect 2167 544 2172 549
rect 2282 558 2287 563
rect 2220 553 2225 558
rect 2188 533 2193 538
rect 2448 601 2453 606
rect 2331 578 2336 583
rect 2332 569 2337 574
rect 2370 544 2375 549
rect 2115 396 2120 401
rect 2150 337 2155 342
rect 2063 323 2068 328
rect 2206 354 2211 359
rect 2206 327 2211 332
rect 2183 321 2188 326
rect 2206 295 2212 300
rect 2164 265 2169 270
rect 2279 279 2284 284
rect 2217 274 2222 279
rect 2185 254 2190 259
rect 2398 322 2403 327
rect 2328 299 2333 304
rect 2329 290 2334 295
rect 2376 265 2381 270
rect 3232 464 3237 469
rect 3247 464 3252 469
rect 3262 464 3267 469
rect 3276 464 3281 469
rect 3247 355 3252 360
rect 3262 348 3267 353
rect 2443 322 2448 327
rect 3248 321 3253 326
rect 2067 62 2072 67
rect 2118 111 2123 116
rect 2153 52 2158 57
rect 2209 69 2214 74
rect 2209 42 2214 47
rect 2186 36 2191 41
rect 2209 10 2215 15
rect 2167 -20 2172 -15
rect 2282 -6 2287 -1
rect 2220 -11 2225 -6
rect 2188 -31 2193 -26
rect 2873 116 2878 121
rect 2919 154 2924 159
rect 2980 155 2985 160
rect 2331 14 2336 19
rect 2332 5 2337 10
rect 2376 -20 2381 -15
rect 1238 -103 1243 -98
rect 455 -139 460 -134
rect 86 -188 92 -182
rect 104 -186 109 -181
rect 363 -184 369 -178
rect 189 -205 195 -200
rect 439 -183 444 -178
rect 395 -205 400 -200
rect 437 -208 442 -203
rect 526 -160 531 -155
rect 504 -168 509 -163
rect 683 -165 688 -160
rect 486 -183 491 -178
rect 449 -225 454 -220
rect 441 -249 446 -244
rect 395 -271 400 -266
rect 820 -165 826 -160
rect 965 -165 971 -160
rect 1090 -165 1095 -160
rect 1315 -165 1320 -160
rect 1374 -160 1379 -155
rect 1524 -160 1529 -155
rect 1663 -160 1668 -155
rect 1787 -160 1792 -155
rect 1462 -165 1467 -160
rect 1601 -165 1606 -160
rect 1725 -165 1730 -160
rect 1238 -187 1243 -182
rect 534 -193 539 -188
rect 485 -249 490 -244
rect 440 -315 445 -310
rect 395 -337 400 -332
rect 2875 -45 2880 -40
rect 2921 -7 2926 -2
rect 2982 -6 2987 -1
rect 3149 43 3154 48
rect 3247 -58 3252 -53
rect 678 -298 683 -293
rect 485 -315 490 -310
rect 815 -298 821 -293
rect 105 -403 110 -398
rect 594 -319 599 -314
rect 960 -298 965 -293
rect 1084 -298 1089 -293
rect 1309 -298 1314 -293
rect 1457 -298 1462 -293
rect 1596 -298 1601 -293
rect 1720 -298 1725 -293
rect 2777 -379 2782 -374
rect 673 -437 678 -432
rect 811 -437 816 -432
rect 873 -433 878 -428
rect 1019 -432 1024 -427
rect 956 -437 961 -432
rect 1080 -437 1085 -432
rect 1143 -433 1148 -428
rect 1305 -437 1310 -432
rect 1453 -437 1458 -432
rect 1592 -437 1597 -432
rect 1716 -437 1721 -432
rect 1833 -481 1838 -476
rect 1834 -586 1839 -581
rect 3262 -78 3267 -73
rect 2892 -122 2897 -117
rect 2874 -199 2879 -194
rect 2920 -161 2925 -156
rect 2981 -160 2986 -155
rect 3276 -160 3281 -155
rect 2874 -347 2879 -342
rect 2920 -309 2925 -304
rect 2981 -308 2986 -303
rect 3416 -347 3421 -342
rect 3386 -405 3391 -400
rect 2927 -435 2932 -430
rect 2927 -502 2932 -497
rect 3144 -506 3149 -501
rect 3462 -431 3467 -426
rect 3335 -511 3340 -506
rect 3345 -511 3350 -506
rect 2856 -567 2861 -562
rect 2919 -569 2924 -564
rect 3120 -583 3125 -578
rect 3319 -525 3324 -520
rect 3491 -430 3496 -425
rect 3195 -586 3200 -581
rect 2898 -636 2903 -631
rect 1834 -708 1839 -703
<< metal2 >>
rect 2125 953 2204 956
rect 2200 914 2204 953
rect 2200 911 2211 914
rect 2160 893 2190 897
rect 1457 877 2067 881
rect 1457 55 1460 877
rect 2186 881 2190 893
rect 2186 876 2188 881
rect 2186 824 2190 876
rect 2200 833 2204 911
rect 2216 911 2217 914
rect 2212 855 2216 882
rect 2303 854 2333 858
rect 2283 834 2284 838
rect 2303 838 2306 854
rect 2289 834 2306 838
rect 2200 829 2222 833
rect 2174 820 2190 824
rect 2334 812 2338 845
rect 2195 809 2338 812
rect 2123 677 2202 680
rect 2198 638 2202 677
rect 2198 635 2209 638
rect 2158 617 2188 621
rect 2184 605 2188 617
rect 1605 598 2067 601
rect 1605 52 1609 598
rect 2184 600 2186 605
rect 2184 548 2188 600
rect 2198 557 2202 635
rect 2214 635 2215 638
rect 2210 579 2214 606
rect 2301 578 2331 582
rect 2281 558 2282 562
rect 2301 562 2304 578
rect 2287 558 2304 562
rect 2198 553 2220 557
rect 2172 544 2188 548
rect 2332 536 2336 569
rect 2371 549 2374 820
rect 2193 533 2336 536
rect 2120 398 2199 401
rect 2195 359 2199 398
rect 2195 356 2206 359
rect 2155 338 2185 342
rect 1757 323 2063 327
rect 2181 326 2185 338
rect 1757 52 1761 323
rect 2181 321 2183 326
rect 2181 269 2185 321
rect 2195 278 2199 356
rect 2211 356 2212 359
rect 2207 300 2211 327
rect 2298 299 2328 303
rect 2278 279 2279 283
rect 2298 283 2301 299
rect 2284 279 2301 283
rect 2195 274 2217 278
rect 2169 265 2185 269
rect 2329 257 2333 290
rect 2370 274 2375 544
rect 2403 324 2443 327
rect 2448 323 2452 601
rect 3233 459 3237 464
rect 3248 459 3252 464
rect 3263 462 3267 464
rect 3277 462 3281 464
rect 2372 271 2379 274
rect 2190 254 2333 257
rect 2376 270 2379 271
rect 2123 113 2202 116
rect 2198 74 2202 113
rect 2198 71 2209 74
rect 1908 63 2067 66
rect 1908 51 1911 63
rect 2158 53 2188 57
rect 2184 41 2188 53
rect 2184 36 2186 41
rect 1403 -15 1411 -12
rect 104 -133 109 -132
rect 86 -182 92 -137
rect 96 -136 109 -133
rect 96 -184 100 -136
rect 137 -141 141 -74
rect 319 -100 366 -97
rect 126 -146 141 -141
rect 252 -116 254 -111
rect 96 -186 104 -184
rect 96 -192 111 -186
rect 104 -398 111 -192
rect 189 -305 195 -205
rect 252 -236 260 -116
rect 319 -178 324 -100
rect 390 -139 394 -132
rect 347 -143 394 -139
rect 455 -142 460 -139
rect 362 -171 369 -143
rect 455 -146 514 -142
rect 509 -155 514 -146
rect 509 -159 526 -155
rect 645 -165 683 -160
rect 787 -165 820 -160
rect 932 -165 965 -160
rect 1058 -165 1090 -160
rect 362 -174 396 -171
rect 319 -181 363 -178
rect 390 -200 396 -174
rect 444 -182 486 -178
rect 390 -205 395 -200
rect 504 -203 508 -168
rect 442 -207 508 -203
rect 523 -191 534 -188
rect 523 -220 527 -191
rect 454 -223 527 -220
rect 252 -240 396 -236
rect 390 -266 396 -240
rect 446 -248 485 -244
rect 390 -271 395 -266
rect 189 -308 396 -305
rect 390 -332 396 -308
rect 445 -314 485 -310
rect 523 -314 527 -223
rect 645 -294 649 -165
rect 645 -298 678 -294
rect 787 -294 791 -165
rect 787 -298 815 -294
rect 932 -294 936 -165
rect 932 -298 960 -294
rect 1058 -294 1062 -165
rect 1239 -182 1243 -103
rect 1403 -156 1407 -15
rect 1545 -17 1558 -14
rect 1379 -160 1407 -156
rect 1523 -160 1524 -156
rect 1545 -156 1549 -17
rect 1683 -18 1709 -15
rect 1529 -160 1549 -156
rect 1683 -156 1686 -18
rect 1714 -18 1715 -15
rect 1842 -19 1861 -16
rect 1668 -160 1686 -156
rect 1786 -160 1787 -156
rect 1842 -156 1846 -19
rect 2184 -16 2188 36
rect 2198 -7 2202 71
rect 2214 71 2215 74
rect 2210 15 2214 42
rect 2301 14 2331 18
rect 2281 -6 2282 -2
rect 2301 -2 2304 14
rect 2287 -6 2304 -2
rect 2198 -11 2220 -7
rect 2172 -20 2188 -16
rect 2332 -28 2336 5
rect 2376 -15 2380 265
rect 2857 199 3175 202
rect 2857 121 2862 199
rect 2924 155 2980 159
rect 2985 155 2986 159
rect 2830 118 2873 121
rect 2193 -31 2336 -28
rect 1792 -160 1846 -156
rect 1277 -165 1315 -160
rect 1428 -165 1462 -160
rect 1566 -165 1601 -160
rect 1695 -165 1725 -160
rect 1058 -298 1084 -294
rect 1277 -294 1281 -165
rect 1277 -298 1309 -294
rect 1428 -294 1432 -165
rect 1428 -298 1457 -294
rect 1566 -294 1570 -165
rect 1566 -298 1596 -294
rect 1695 -294 1699 -165
rect 1695 -298 1720 -294
rect 523 -318 594 -314
rect 390 -337 395 -332
rect 104 -402 105 -398
rect 110 -402 111 -398
rect 645 -433 649 -298
rect 645 -437 673 -433
rect 787 -433 791 -298
rect 871 -432 873 -428
rect 787 -437 811 -433
rect 878 -432 888 -428
rect 884 -703 888 -432
rect 932 -433 936 -298
rect 1018 -432 1019 -428
rect 1024 -432 1031 -428
rect 932 -437 956 -433
rect 1028 -581 1031 -432
rect 1058 -433 1062 -298
rect 1142 -432 1143 -428
rect 1058 -437 1080 -433
rect 1148 -432 1157 -428
rect 1154 -476 1157 -432
rect 1277 -433 1281 -298
rect 1277 -437 1305 -433
rect 1428 -433 1432 -298
rect 1428 -437 1453 -433
rect 1566 -433 1570 -298
rect 1566 -437 1592 -433
rect 1695 -433 1699 -298
rect 2830 -375 2833 118
rect 2859 45 3149 48
rect 2859 -40 2862 45
rect 2926 -6 2982 -2
rect 2987 -6 2988 -2
rect 2782 -378 2833 -375
rect 1695 -437 1716 -433
rect 1154 -481 1833 -476
rect 1028 -586 1834 -581
rect 2830 -631 2833 -378
rect 2847 -43 2875 -40
rect 2847 -564 2850 -43
rect 2857 -121 2892 -117
rect 2857 -194 2860 -121
rect 2925 -160 2981 -156
rect 2986 -160 2987 -156
rect 2857 -197 2874 -194
rect 2857 -496 2860 -197
rect 3233 -269 3236 459
rect 3248 360 3251 459
rect 3248 326 3251 355
rect 3263 353 3266 462
rect 3248 -53 3251 321
rect 2865 -272 3236 -269
rect 2865 -342 2868 -272
rect 2925 -308 2981 -304
rect 2986 -308 2987 -304
rect 2865 -345 2874 -342
rect 2865 -431 2868 -345
rect 2865 -435 2927 -431
rect 2861 -501 2927 -497
rect 3120 -504 3144 -501
rect 2847 -567 2856 -564
rect 2861 -567 2919 -564
rect 2847 -568 2919 -567
rect 3120 -578 3124 -504
rect 3248 -564 3251 -58
rect 3263 -73 3266 348
rect 3263 -520 3266 -78
rect 3277 -155 3280 462
rect 3277 -415 3280 -160
rect 3387 -345 3416 -342
rect 3387 -400 3390 -345
rect 3277 -418 3418 -415
rect 3415 -426 3418 -418
rect 3415 -429 3462 -426
rect 3336 -520 3340 -511
rect 3263 -523 3319 -520
rect 3324 -523 3340 -520
rect 3346 -564 3350 -511
rect 3492 -564 3496 -430
rect 3248 -567 3496 -564
rect 3248 -581 3251 -567
rect 3200 -584 3251 -581
rect 2830 -635 2898 -631
rect 884 -708 1834 -703
<< m3contact >>
rect 3175 197 3180 202
<< m123contact >>
rect 2077 862 2082 867
rect 2075 584 2080 589
rect 2072 308 2077 313
rect 2973 485 2978 490
rect 2981 442 2986 447
rect 2972 419 2977 424
rect 2981 376 2986 381
rect 2972 352 2977 357
rect 2981 309 2986 314
rect 2972 285 2977 290
rect 2075 32 2080 37
rect 1482 -9 1487 -4
rect 1631 -11 1636 -6
rect 744 -160 749 -155
rect 882 -161 887 -155
rect 1028 -161 1033 -156
rect 1152 -161 1157 -156
rect 1783 -12 1788 -7
rect 1933 -13 1938 -8
rect 2120 -21 2125 -16
rect 2981 242 2986 247
rect 2972 179 2977 184
rect 1852 -186 1857 -181
rect 2762 -351 2767 -346
rect 2981 96 2986 101
rect 2972 18 2977 23
rect 3007 18 3012 23
rect 2982 -24 2987 -19
rect 2751 -540 2757 -535
rect 2972 -136 2977 -131
rect 2981 -178 2986 -173
rect 2972 -284 2977 -279
rect 2981 -326 2986 -321
rect 2972 -410 2977 -405
rect 2981 -453 2986 -448
rect 2972 -476 2977 -471
rect 2856 -501 2861 -496
rect 2981 -519 2986 -514
rect 2868 -530 2874 -524
rect 2972 -543 2977 -538
rect 3233 -506 3238 -501
rect 3234 -539 3239 -534
rect 3633 295 3638 300
rect 3580 -32 3585 -27
rect 3658 -94 3663 -89
rect 3684 -358 3689 -353
rect 3285 -431 3290 -426
rect 2981 -586 2986 -581
rect 2972 -610 2977 -605
rect 2981 -653 2986 -648
<< metal3 >>
rect 759 862 2077 867
rect 759 859 2079 862
rect 742 -160 744 -156
rect 759 -156 768 859
rect 893 589 902 590
rect 1040 589 1049 590
rect 1172 589 1181 590
rect 893 586 2075 589
rect 749 -160 768 -156
rect 881 -160 882 -156
rect 893 -156 902 586
rect 2973 424 2977 485
rect 2973 357 2977 419
rect 1040 309 2072 313
rect 1040 -156 1049 309
rect 2973 290 2977 352
rect 2973 184 2977 285
rect 1172 111 1181 134
rect 1172 104 2043 111
rect 1172 -156 1181 104
rect 2035 38 2043 104
rect 2035 37 2078 38
rect 2035 35 2075 37
rect 2973 23 2977 179
rect 1483 -55 1486 -9
rect 1632 -55 1636 -11
rect 1784 -55 1788 -12
rect 1934 -31 1937 -13
rect 2115 -21 2120 -18
rect 2115 -31 2118 -21
rect 1934 -34 2118 -31
rect 1934 -55 1937 -34
rect 1483 -58 1937 -55
rect 887 -160 902 -156
rect 1027 -160 1028 -156
rect 1033 -160 1049 -156
rect 1151 -160 1152 -156
rect 1157 -160 1181 -156
rect 1853 -181 1856 -58
rect 2973 -131 2977 18
rect 2973 -279 2977 -136
rect 2767 -350 2872 -346
rect 2869 -490 2872 -350
rect 2973 -405 2977 -284
rect 2973 -471 2977 -410
rect 2857 -536 2860 -501
rect 2869 -524 2873 -490
rect 2757 -539 2860 -536
rect 2973 -538 2977 -476
rect 2973 -605 2977 -543
rect 2981 381 2985 442
rect 2981 314 2985 376
rect 2981 247 2985 309
rect 2981 101 2985 242
rect 3634 202 3638 295
rect 3180 198 3638 202
rect 2981 -19 2985 96
rect 3012 19 3580 23
rect 2981 -24 2982 -19
rect 2981 -173 2985 -24
rect 3576 -30 3580 19
rect 2981 -191 2985 -178
rect 3659 -191 3663 -94
rect 2981 -194 3663 -191
rect 2981 -321 2985 -194
rect 2981 -448 2985 -326
rect 3234 -429 3285 -426
rect 2981 -514 2985 -453
rect 3234 -501 3237 -429
rect 2981 -581 2985 -519
rect 3685 -534 3689 -358
rect 3239 -538 3689 -534
rect 2981 -648 2985 -586
<< labels >>
rlabel metal1 97 -72 98 -71 1 VDD
rlabel metal1 88 -114 89 -113 1 s0
rlabel metal1 80 -169 81 -168 1 s1
rlabel metal1 90 -404 91 -403 1 gnd
rlabel m2contact 439 -206 440 -205 1 d1
rlabel metal1 439 -271 440 -270 1 d2
rlabel metal1 439 -337 440 -336 1 d3
rlabel metal1 438 -136 439 -135 1 d0
rlabel metal1 688 -163 688 -163 1 a0
rlabel metal1 826 -163 826 -163 1 a1
rlabel metal1 971 -163 971 -163 1 a2
rlabel metal1 1096 -163 1096 -163 1 a3
rlabel metal1 1320 -163 1320 -163 1 b0
rlabel metal1 1467 -162 1467 -162 1 b1
rlabel metal1 1606 -162 1606 -162 1 b2
rlabel metal1 1730 -162 1730 -162 1 b3
rlabel metal1 881 -158 881 -158 1 ena1as
rlabel metal1 1027 -158 1027 -158 1 ena2as
rlabel metal1 1151 -158 1151 -158 1 ena3as
rlabel m2contact 1376 -158 1376 -158 1 enb0as
rlabel metal1 1662 -158 1662 -158 1 enb2as
rlabel metal1 1786 -158 1786 -158 1 enb3as
rlabel metal1 738 -291 738 -291 1 ena0c
rlabel metal1 877 -291 877 -291 1 ena1c
rlabel metal1 1022 -291 1022 -291 1 ena2c
rlabel metal1 1146 -291 1146 -291 1 ena3c
rlabel metal1 1371 -291 1371 -291 1 enb0c
rlabel metal1 1518 -291 1518 -291 1 enb1c
rlabel metal1 1657 -291 1657 -291 1 enb2c
rlabel metal1 1781 -291 1781 -291 1 enb3c
rlabel metal1 734 -430 734 -430 1 ena0a
rlabel metal1 1018 -430 1018 -430 1 ena2a
rlabel metal1 1142 -430 1142 -430 1 ena3a
rlabel metal1 1367 -430 1367 -430 1 enb0a
rlabel metal1 1514 -430 1514 -430 1 enb1a
rlabel metal1 1653 -430 1653 -430 1 enb2a
rlabel metal1 1777 -430 1777 -430 1 enb3a
rlabel metal1 1893 -808 1893 -808 1 and0
rlabel metal1 1893 -701 1893 -701 1 and1
rlabel metal1 1893 -579 1893 -579 1 and2
rlabel metal1 1893 -474 1893 -474 1 and3
rlabel metal1 872 -430 872 -430 1 ena1a
rlabel metal1 1523 -158 1523 -158 1 enb1as
rlabel metal1 743 -158 743 -158 1 ena0as
rlabel metal1 2243 949 2243 950 1 sout0
rlabel metal1 2240 673 2240 674 1 sout1
rlabel metal1 2236 395 2236 396 1 sout2
rlabel metal1 2239 109 2239 110 1 sout3
rlabel metal1 2413 15 2413 15 1 cout
rlabel metal1 3740 467 3740 467 7 gtr
rlabel metal1 3731 -313 3731 -313 1 lsr
rlabel polysilicon 3660 -341 3660 -341 1 w1
rlabel polysilicon 3672 -341 3672 -341 1 w2
rlabel polysilicon 3687 -341 3687 -341 1 w3
rlabel polysilicon 3697 -341 3697 -341 1 w4
rlabel metal1 3775 -59 3775 -59 1 equ
rlabel metal1 3697 -61 3697 -61 1 pequ
rlabel metal1 3177 -582 3177 -582 1 check1
rlabel metal1 3016 157 3016 157 1 x3
rlabel metal1 3018 -4 3018 -4 1 x2
rlabel metal1 3018 -158 3018 -158 1 x1
rlabel metal1 3016 -306 3016 -306 1 x0
<< end >>
